// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jul 13 2021 16:01:58

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    PORT1,
    CLK,
    BUT2,
    BUT1);

    output PORT1;
    input CLK;
    input BUT2;
    input BUT1;

    wire N__2680;
    wire N__2679;
    wire N__2678;
    wire N__2669;
    wire N__2668;
    wire N__2667;
    wire N__2660;
    wire N__2659;
    wire N__2658;
    wire N__2651;
    wire N__2650;
    wire N__2649;
    wire N__2632;
    wire N__2631;
    wire N__2628;
    wire N__2627;
    wire N__2626;
    wire N__2619;
    wire N__2616;
    wire N__2613;
    wire N__2610;
    wire N__2607;
    wire N__2604;
    wire N__2601;
    wire N__2598;
    wire N__2593;
    wire N__2592;
    wire N__2589;
    wire N__2586;
    wire N__2583;
    wire N__2580;
    wire N__2575;
    wire N__2574;
    wire N__2573;
    wire N__2570;
    wire N__2565;
    wire N__2560;
    wire N__2559;
    wire N__2558;
    wire N__2555;
    wire N__2550;
    wire N__2547;
    wire N__2542;
    wire N__2541;
    wire N__2540;
    wire N__2539;
    wire N__2536;
    wire N__2531;
    wire N__2528;
    wire N__2521;
    wire N__2520;
    wire N__2519;
    wire N__2518;
    wire N__2515;
    wire N__2508;
    wire N__2503;
    wire N__2500;
    wire N__2499;
    wire N__2496;
    wire N__2493;
    wire N__2492;
    wire N__2491;
    wire N__2488;
    wire N__2485;
    wire N__2480;
    wire N__2473;
    wire N__2470;
    wire N__2467;
    wire N__2466;
    wire N__2463;
    wire N__2460;
    wire N__2455;
    wire N__2452;
    wire N__2449;
    wire N__2446;
    wire N__2443;
    wire N__2440;
    wire N__2439;
    wire N__2436;
    wire N__2433;
    wire N__2428;
    wire N__2427;
    wire N__2424;
    wire N__2423;
    wire N__2420;
    wire N__2415;
    wire N__2410;
    wire N__2409;
    wire N__2406;
    wire N__2405;
    wire N__2402;
    wire N__2401;
    wire N__2398;
    wire N__2391;
    wire N__2386;
    wire N__2383;
    wire N__2380;
    wire N__2377;
    wire N__2376;
    wire N__2371;
    wire N__2370;
    wire N__2369;
    wire N__2366;
    wire N__2363;
    wire N__2362;
    wire N__2361;
    wire N__2358;
    wire N__2355;
    wire N__2352;
    wire N__2347;
    wire N__2344;
    wire N__2335;
    wire N__2334;
    wire N__2331;
    wire N__2330;
    wire N__2327;
    wire N__2326;
    wire N__2325;
    wire N__2322;
    wire N__2319;
    wire N__2316;
    wire N__2313;
    wire N__2310;
    wire N__2309;
    wire N__2306;
    wire N__2303;
    wire N__2298;
    wire N__2295;
    wire N__2292;
    wire N__2289;
    wire N__2286;
    wire N__2281;
    wire N__2278;
    wire N__2269;
    wire N__2266;
    wire N__2263;
    wire N__2262;
    wire N__2261;
    wire N__2260;
    wire N__2257;
    wire N__2250;
    wire N__2245;
    wire N__2244;
    wire N__2241;
    wire N__2238;
    wire N__2235;
    wire N__2230;
    wire N__2227;
    wire N__2226;
    wire N__2223;
    wire N__2220;
    wire N__2217;
    wire N__2212;
    wire N__2209;
    wire N__2206;
    wire N__2205;
    wire N__2202;
    wire N__2199;
    wire N__2194;
    wire N__2193;
    wire N__2192;
    wire N__2191;
    wire N__2190;
    wire N__2189;
    wire N__2188;
    wire N__2187;
    wire N__2186;
    wire N__2185;
    wire N__2184;
    wire N__2161;
    wire N__2158;
    wire N__2155;
    wire N__2152;
    wire N__2149;
    wire N__2148;
    wire N__2145;
    wire N__2142;
    wire N__2137;
    wire N__2134;
    wire N__2133;
    wire N__2130;
    wire N__2127;
    wire N__2126;
    wire N__2125;
    wire N__2120;
    wire N__2115;
    wire N__2110;
    wire N__2107;
    wire N__2104;
    wire N__2101;
    wire N__2098;
    wire N__2097;
    wire N__2096;
    wire N__2095;
    wire N__2092;
    wire N__2087;
    wire N__2084;
    wire N__2079;
    wire N__2074;
    wire N__2073;
    wire N__2072;
    wire N__2071;
    wire N__2068;
    wire N__2063;
    wire N__2060;
    wire N__2053;
    wire N__2052;
    wire N__2051;
    wire N__2048;
    wire N__2045;
    wire N__2042;
    wire N__2035;
    wire N__2034;
    wire N__2033;
    wire N__2032;
    wire N__2029;
    wire N__2026;
    wire N__2023;
    wire N__2020;
    wire N__2017;
    wire N__2014;
    wire N__2005;
    wire N__2004;
    wire N__2001;
    wire N__1998;
    wire N__1995;
    wire N__1990;
    wire N__1987;
    wire N__1986;
    wire N__1983;
    wire N__1980;
    wire N__1977;
    wire N__1972;
    wire N__1969;
    wire N__1968;
    wire N__1965;
    wire N__1962;
    wire N__1959;
    wire N__1954;
    wire N__1951;
    wire N__1950;
    wire N__1947;
    wire N__1944;
    wire N__1941;
    wire N__1936;
    wire N__1933;
    wire N__1932;
    wire N__1929;
    wire N__1926;
    wire N__1923;
    wire N__1918;
    wire N__1915;
    wire N__1914;
    wire N__1911;
    wire N__1908;
    wire N__1905;
    wire N__1900;
    wire N__1897;
    wire N__1894;
    wire N__1893;
    wire N__1890;
    wire N__1887;
    wire N__1882;
    wire N__1879;
    wire N__1876;
    wire N__1873;
    wire N__1870;
    wire N__1869;
    wire N__1866;
    wire N__1863;
    wire N__1858;
    wire N__1855;
    wire N__1852;
    wire N__1851;
    wire N__1850;
    wire N__1849;
    wire N__1846;
    wire N__1843;
    wire N__1840;
    wire N__1837;
    wire N__1836;
    wire N__1833;
    wire N__1828;
    wire N__1825;
    wire N__1822;
    wire N__1813;
    wire N__1810;
    wire N__1809;
    wire N__1808;
    wire N__1805;
    wire N__1802;
    wire N__1799;
    wire N__1794;
    wire N__1793;
    wire N__1792;
    wire N__1791;
    wire N__1790;
    wire N__1789;
    wire N__1786;
    wire N__1783;
    wire N__1774;
    wire N__1771;
    wire N__1762;
    wire N__1761;
    wire N__1758;
    wire N__1757;
    wire N__1756;
    wire N__1753;
    wire N__1750;
    wire N__1745;
    wire N__1738;
    wire N__1737;
    wire N__1736;
    wire N__1735;
    wire N__1732;
    wire N__1729;
    wire N__1726;
    wire N__1723;
    wire N__1714;
    wire N__1713;
    wire N__1712;
    wire N__1711;
    wire N__1710;
    wire N__1707;
    wire N__1702;
    wire N__1699;
    wire N__1696;
    wire N__1687;
    wire N__1686;
    wire N__1685;
    wire N__1682;
    wire N__1677;
    wire N__1672;
    wire N__1671;
    wire N__1670;
    wire N__1669;
    wire N__1668;
    wire N__1665;
    wire N__1662;
    wire N__1661;
    wire N__1660;
    wire N__1657;
    wire N__1654;
    wire N__1651;
    wire N__1648;
    wire N__1643;
    wire N__1638;
    wire N__1635;
    wire N__1624;
    wire N__1623;
    wire N__1620;
    wire N__1617;
    wire N__1612;
    wire N__1609;
    wire N__1606;
    wire N__1603;
    wire N__1602;
    wire N__1601;
    wire N__1600;
    wire N__1597;
    wire N__1594;
    wire N__1591;
    wire N__1588;
    wire N__1585;
    wire N__1576;
    wire N__1573;
    wire N__1572;
    wire N__1569;
    wire N__1566;
    wire N__1561;
    wire N__1560;
    wire N__1557;
    wire N__1556;
    wire N__1553;
    wire N__1550;
    wire N__1545;
    wire N__1540;
    wire N__1537;
    wire N__1534;
    wire N__1533;
    wire N__1532;
    wire N__1529;
    wire N__1526;
    wire N__1523;
    wire N__1516;
    wire N__1513;
    wire N__1510;
    wire N__1507;
    wire N__1504;
    wire N__1503;
    wire N__1498;
    wire N__1495;
    wire N__1492;
    wire N__1489;
    wire N__1486;
    wire N__1485;
    wire N__1484;
    wire N__1483;
    wire N__1482;
    wire N__1473;
    wire N__1470;
    wire N__1465;
    wire N__1464;
    wire N__1463;
    wire N__1462;
    wire N__1461;
    wire N__1460;
    wire N__1449;
    wire N__1446;
    wire N__1441;
    wire N__1440;
    wire N__1439;
    wire N__1438;
    wire N__1437;
    wire N__1428;
    wire N__1425;
    wire N__1420;
    wire N__1417;
    wire N__1414;
    wire N__1411;
    wire N__1408;
    wire N__1407;
    wire N__1402;
    wire N__1399;
    wire N__1396;
    wire N__1393;
    wire N__1390;
    wire N__1389;
    wire N__1386;
    wire N__1383;
    wire N__1378;
    wire N__1375;
    wire N__1374;
    wire N__1371;
    wire N__1368;
    wire N__1363;
    wire N__1362;
    wire N__1359;
    wire N__1356;
    wire N__1351;
    wire N__1350;
    wire N__1347;
    wire N__1344;
    wire N__1339;
    wire N__1338;
    wire N__1335;
    wire N__1332;
    wire N__1327;
    wire N__1324;
    wire N__1323;
    wire N__1320;
    wire N__1317;
    wire N__1312;
    wire N__1311;
    wire N__1308;
    wire N__1305;
    wire N__1300;
    wire N__1297;
    wire N__1294;
    wire N__1291;
    wire N__1288;
    wire N__1285;
    wire N__1282;
    wire N__1279;
    wire N__1276;
    wire N__1273;
    wire N__1270;
    wire N__1269;
    wire N__1266;
    wire N__1263;
    wire N__1258;
    wire N__1257;
    wire N__1254;
    wire N__1251;
    wire N__1246;
    wire N__1245;
    wire N__1242;
    wire N__1239;
    wire N__1234;
    wire N__1233;
    wire N__1230;
    wire N__1227;
    wire N__1222;
    wire N__1219;
    wire N__1216;
    wire N__1213;
    wire N__1210;
    wire N__1207;
    wire N__1204;
    wire N__1201;
    wire N__1200;
    wire N__1195;
    wire N__1192;
    wire N__1191;
    wire N__1186;
    wire N__1183;
    wire N__1180;
    wire N__1179;
    wire N__1174;
    wire N__1171;
    wire N__1170;
    wire N__1165;
    wire N__1162;
    wire N__1159;
    wire N__1156;
    wire N__1153;
    wire N__1150;
    wire N__1147;
    wire N__1144;
    wire N__1141;
    wire GNDG0;
    wire VCCG0;
    wire bfn_1_2_0_;
    wire delay_cry_0;
    wire delay_cry_1;
    wire delay_cry_2;
    wire delay_cry_3;
    wire delay_cry_4;
    wire delay_cry_5;
    wire delay_cry_6;
    wire delay_cry_7;
    wire bfn_1_3_0_;
    wire delay_cry_8;
    wire delay_cry_9;
    wire delay_cry_10;
    wire delay_cry_11;
    wire delay_cry_12;
    wire delay_cry_13;
    wire delayZ0Z_14;
    wire delayZ0Z_13;
    wire delayZ0Z_12;
    wire delayZ0Z_11;
    wire bfn_1_7_0_;
    wire clk_div_2_cry_1;
    wire clk_div_2_cry_2;
    wire clk_div_2_cry_3;
    wire clk_div_2_cry_4;
    wire clk_div_2_cry_5;
    wire clk_div_2_cry_6;
    wire clk_div_2_cry_7;
    wire clk_div_2_cry_8;
    wire bfn_1_8_0_;
    wire clk_div_2_cry_9;
    wire clk_div_2_cry_10;
    wire delayZ0Z_6;
    wire delayZ0Z_5;
    wire delayZ0Z_4;
    wire delayZ0Z_7;
    wire delayZ0Z_10;
    wire delayZ0Z_8;
    wire delayZ0Z_9;
    wire delayZ0Z_0;
    wire delayZ0Z_3;
    wire delayZ0Z_1;
    wire delayZ0Z_2;
    wire un1_ten_ms_7;
    wire un1_ten_ms_9;
    wire un1_ten_ms_8_cascade_;
    wire un1_ten_ms_10;
    wire how_1_c2;
    wire PWM_NUMZ0Z_3;
    wire PWM_NUMZ0Z_1;
    wire howZ0Z_0;
    wire howZ0Z_2;
    wire howZ0Z_1;
    wire PWM_NUMZ0Z_2;
    wire PORT_r3_2;
    wire PORT_r3_3;
    wire g0_2;
    wire g0_4_cascade_;
    wire PWM_NUM_RNIKTNT2Z0Z_0;
    wire PWM_NUM_RNIKTNT2Z0Z_0_cascade_;
    wire N_78_0;
    wire PWM_NUMZ0Z_4;
    wire g0_3;
    wire cntrZ0Z_4;
    wire clk_div_RNIM1KP1Z0Z_11;
    wire cntrZ0Z_3;
    wire cntrZ0Z_2;
    wire cntrZ0Z_1;
    wire un2_cntr_c4;
    wire cntrZ0Z_0;
    wire PWM_NUMZ0Z_0;
    wire un1_cntr_0;
    wire cntrZ0Z_5;
    wire PWM_NUMZ0Z_5;
    wire cntrZ0Z_6;
    wire PORT1_c;
    wire PORT_r3_1;
    wire clk_div_RNI06L91Z0Z_11;
    wire clk_div_i_11;
    wire clk_divZ0Z_1;
    wire clk_divZ0Z_0;
    wire bfn_2_8_0_;
    wire clk_divZ0Z_2;
    wire clk_div_1_cry_1;
    wire clk_divZ0Z_3;
    wire clk_div_1_cry_2;
    wire clk_divZ0Z_4;
    wire clk_div_1_cry_3;
    wire clk_divZ0Z_5;
    wire clk_div_1_cry_4;
    wire clk_divZ0Z_6;
    wire clk_div_1_cry_5;
    wire clk_divZ0Z_7;
    wire clk_div_1_cry_6;
    wire clk_divZ0Z_8;
    wire clk_div_1_cry_7;
    wire clk_div_1_cry_8;
    wire clk_divZ0Z_9;
    wire bfn_2_9_0_;
    wire clk_div_1_cry_9;
    wire clk_divZ0Z_10;
    wire CLK_0_c_g;
    wire upZ0Z_2;
    wire upZ0Z_1;
    wire shift_ret_1_RNI69IQZ0;
    wire BUT1_c;
    wire level_0;
    wire shift_0Z0Z_1;
    wire upZ0Z_0;
    wire shift_0Z0Z_2;
    wire downZ0Z_1;
    wire downZ0Z_2;
    wire shift2_ret_1_RNITCIZ0Z51;
    wire level2_0;
    wire shift2_0Z0Z_1;
    wire BUT2_c;
    wire downZ0Z_0;
    wire un1_ten_ms_i;
    wire shift2_0Z0Z_2;
    wire _gnd_net_;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__2678),
            .GLOBALBUFFEROUTPUT(CLK_0_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__2680),
            .DIN(N__2679),
            .DOUT(N__2678),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__2680),
            .PADOUT(N__2679),
            .PADIN(N__2678),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PORT1_obuf_iopad (
            .OE(N__2669),
            .DIN(N__2668),
            .DOUT(N__2667),
            .PACKAGEPIN(PORT1));
    defparam PORT1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PORT1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PORT1_obuf_preio (
            .PADOEN(N__2669),
            .PADOUT(N__2668),
            .PADIN(N__2667),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1540),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUT2_ibuf_iopad (
            .OE(N__2660),
            .DIN(N__2659),
            .DOUT(N__2658),
            .PACKAGEPIN(BUT2));
    defparam BUT2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BUT2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BUT2_ibuf_preio (
            .PADOEN(N__2660),
            .PADOUT(N__2659),
            .PADIN(N__2658),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BUT2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUT1_ibuf_iopad (
            .OE(N__2651),
            .DIN(N__2650),
            .DOUT(N__2649),
            .PACKAGEPIN(BUT1));
    defparam BUT1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BUT1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BUT1_ibuf_preio (
            .PADOEN(N__2651),
            .PADOUT(N__2650),
            .PADIN(N__2649),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BUT1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__597 (
            .O(N__2632),
            .I(N__2628));
    InMux I__596 (
            .O(N__2631),
            .I(N__2619));
    InMux I__595 (
            .O(N__2628),
            .I(N__2619));
    InMux I__594 (
            .O(N__2627),
            .I(N__2619));
    InMux I__593 (
            .O(N__2626),
            .I(N__2616));
    LocalMux I__592 (
            .O(N__2619),
            .I(N__2613));
    LocalMux I__591 (
            .O(N__2616),
            .I(N__2610));
    Span4Mux_h I__590 (
            .O(N__2613),
            .I(N__2607));
    Span4Mux_v I__589 (
            .O(N__2610),
            .I(N__2604));
    Span4Mux_h I__588 (
            .O(N__2607),
            .I(N__2601));
    Span4Mux_h I__587 (
            .O(N__2604),
            .I(N__2598));
    Odrv4 I__586 (
            .O(N__2601),
            .I(BUT1_c));
    Odrv4 I__585 (
            .O(N__2598),
            .I(BUT1_c));
    CascadeMux I__584 (
            .O(N__2593),
            .I(N__2589));
    CascadeMux I__583 (
            .O(N__2592),
            .I(N__2586));
    InMux I__582 (
            .O(N__2589),
            .I(N__2583));
    InMux I__581 (
            .O(N__2586),
            .I(N__2580));
    LocalMux I__580 (
            .O(N__2583),
            .I(level_0));
    LocalMux I__579 (
            .O(N__2580),
            .I(level_0));
    InMux I__578 (
            .O(N__2575),
            .I(N__2570));
    InMux I__577 (
            .O(N__2574),
            .I(N__2565));
    InMux I__576 (
            .O(N__2573),
            .I(N__2565));
    LocalMux I__575 (
            .O(N__2570),
            .I(shift_0Z0Z_1));
    LocalMux I__574 (
            .O(N__2565),
            .I(shift_0Z0Z_1));
    CascadeMux I__573 (
            .O(N__2560),
            .I(N__2555));
    InMux I__572 (
            .O(N__2559),
            .I(N__2550));
    InMux I__571 (
            .O(N__2558),
            .I(N__2550));
    InMux I__570 (
            .O(N__2555),
            .I(N__2547));
    LocalMux I__569 (
            .O(N__2550),
            .I(N__2542));
    LocalMux I__568 (
            .O(N__2547),
            .I(N__2542));
    Span4Mux_v I__567 (
            .O(N__2542),
            .I(N__2536));
    InMux I__566 (
            .O(N__2541),
            .I(N__2531));
    InMux I__565 (
            .O(N__2540),
            .I(N__2531));
    InMux I__564 (
            .O(N__2539),
            .I(N__2528));
    Odrv4 I__563 (
            .O(N__2536),
            .I(upZ0Z_0));
    LocalMux I__562 (
            .O(N__2531),
            .I(upZ0Z_0));
    LocalMux I__561 (
            .O(N__2528),
            .I(upZ0Z_0));
    CEMux I__560 (
            .O(N__2521),
            .I(N__2515));
    InMux I__559 (
            .O(N__2520),
            .I(N__2508));
    InMux I__558 (
            .O(N__2519),
            .I(N__2508));
    InMux I__557 (
            .O(N__2518),
            .I(N__2508));
    LocalMux I__556 (
            .O(N__2515),
            .I(shift_0Z0Z_2));
    LocalMux I__555 (
            .O(N__2508),
            .I(shift_0Z0Z_2));
    InMux I__554 (
            .O(N__2503),
            .I(N__2500));
    LocalMux I__553 (
            .O(N__2500),
            .I(N__2496));
    InMux I__552 (
            .O(N__2499),
            .I(N__2493));
    Span4Mux_v I__551 (
            .O(N__2496),
            .I(N__2488));
    LocalMux I__550 (
            .O(N__2493),
            .I(N__2485));
    InMux I__549 (
            .O(N__2492),
            .I(N__2480));
    InMux I__548 (
            .O(N__2491),
            .I(N__2480));
    Odrv4 I__547 (
            .O(N__2488),
            .I(downZ0Z_1));
    Odrv12 I__546 (
            .O(N__2485),
            .I(downZ0Z_1));
    LocalMux I__545 (
            .O(N__2480),
            .I(downZ0Z_1));
    InMux I__544 (
            .O(N__2473),
            .I(N__2470));
    LocalMux I__543 (
            .O(N__2470),
            .I(N__2467));
    Span4Mux_v I__542 (
            .O(N__2467),
            .I(N__2463));
    InMux I__541 (
            .O(N__2466),
            .I(N__2460));
    Odrv4 I__540 (
            .O(N__2463),
            .I(downZ0Z_2));
    LocalMux I__539 (
            .O(N__2460),
            .I(downZ0Z_2));
    CEMux I__538 (
            .O(N__2455),
            .I(N__2452));
    LocalMux I__537 (
            .O(N__2452),
            .I(N__2449));
    Span4Mux_v I__536 (
            .O(N__2449),
            .I(N__2446));
    Span4Mux_s0_v I__535 (
            .O(N__2446),
            .I(N__2443));
    Odrv4 I__534 (
            .O(N__2443),
            .I(shift2_ret_1_RNITCIZ0Z51));
    InMux I__533 (
            .O(N__2440),
            .I(N__2436));
    InMux I__532 (
            .O(N__2439),
            .I(N__2433));
    LocalMux I__531 (
            .O(N__2436),
            .I(level2_0));
    LocalMux I__530 (
            .O(N__2433),
            .I(level2_0));
    CascadeMux I__529 (
            .O(N__2428),
            .I(N__2424));
    InMux I__528 (
            .O(N__2427),
            .I(N__2420));
    InMux I__527 (
            .O(N__2424),
            .I(N__2415));
    InMux I__526 (
            .O(N__2423),
            .I(N__2415));
    LocalMux I__525 (
            .O(N__2420),
            .I(shift2_0Z0Z_1));
    LocalMux I__524 (
            .O(N__2415),
            .I(shift2_0Z0Z_1));
    InMux I__523 (
            .O(N__2410),
            .I(N__2406));
    CascadeMux I__522 (
            .O(N__2409),
            .I(N__2402));
    LocalMux I__521 (
            .O(N__2406),
            .I(N__2398));
    InMux I__520 (
            .O(N__2405),
            .I(N__2391));
    InMux I__519 (
            .O(N__2402),
            .I(N__2391));
    InMux I__518 (
            .O(N__2401),
            .I(N__2391));
    Span4Mux_v I__517 (
            .O(N__2398),
            .I(N__2386));
    LocalMux I__516 (
            .O(N__2391),
            .I(N__2386));
    Span4Mux_h I__515 (
            .O(N__2386),
            .I(N__2383));
    Odrv4 I__514 (
            .O(N__2383),
            .I(BUT2_c));
    CascadeMux I__513 (
            .O(N__2380),
            .I(N__2377));
    InMux I__512 (
            .O(N__2377),
            .I(N__2371));
    InMux I__511 (
            .O(N__2376),
            .I(N__2371));
    LocalMux I__510 (
            .O(N__2371),
            .I(N__2366));
    InMux I__509 (
            .O(N__2370),
            .I(N__2363));
    CascadeMux I__508 (
            .O(N__2369),
            .I(N__2358));
    Span4Mux_v I__507 (
            .O(N__2366),
            .I(N__2355));
    LocalMux I__506 (
            .O(N__2363),
            .I(N__2352));
    InMux I__505 (
            .O(N__2362),
            .I(N__2347));
    InMux I__504 (
            .O(N__2361),
            .I(N__2347));
    InMux I__503 (
            .O(N__2358),
            .I(N__2344));
    Odrv4 I__502 (
            .O(N__2355),
            .I(downZ0Z_0));
    Odrv12 I__501 (
            .O(N__2352),
            .I(downZ0Z_0));
    LocalMux I__500 (
            .O(N__2347),
            .I(downZ0Z_0));
    LocalMux I__499 (
            .O(N__2344),
            .I(downZ0Z_0));
    ClkMux I__498 (
            .O(N__2335),
            .I(N__2331));
    ClkMux I__497 (
            .O(N__2334),
            .I(N__2327));
    LocalMux I__496 (
            .O(N__2331),
            .I(N__2322));
    ClkMux I__495 (
            .O(N__2330),
            .I(N__2319));
    LocalMux I__494 (
            .O(N__2327),
            .I(N__2316));
    ClkMux I__493 (
            .O(N__2326),
            .I(N__2313));
    ClkMux I__492 (
            .O(N__2325),
            .I(N__2310));
    Span4Mux_s3_v I__491 (
            .O(N__2322),
            .I(N__2306));
    LocalMux I__490 (
            .O(N__2319),
            .I(N__2303));
    Span4Mux_v I__489 (
            .O(N__2316),
            .I(N__2298));
    LocalMux I__488 (
            .O(N__2313),
            .I(N__2298));
    LocalMux I__487 (
            .O(N__2310),
            .I(N__2295));
    ClkMux I__486 (
            .O(N__2309),
            .I(N__2292));
    Span4Mux_h I__485 (
            .O(N__2306),
            .I(N__2289));
    Span4Mux_v I__484 (
            .O(N__2303),
            .I(N__2286));
    Span4Mux_h I__483 (
            .O(N__2298),
            .I(N__2281));
    Span4Mux_h I__482 (
            .O(N__2295),
            .I(N__2281));
    LocalMux I__481 (
            .O(N__2292),
            .I(N__2278));
    Odrv4 I__480 (
            .O(N__2289),
            .I(un1_ten_ms_i));
    Odrv4 I__479 (
            .O(N__2286),
            .I(un1_ten_ms_i));
    Odrv4 I__478 (
            .O(N__2281),
            .I(un1_ten_ms_i));
    Odrv12 I__477 (
            .O(N__2278),
            .I(un1_ten_ms_i));
    CEMux I__476 (
            .O(N__2269),
            .I(N__2266));
    LocalMux I__475 (
            .O(N__2266),
            .I(N__2263));
    Sp12to4 I__474 (
            .O(N__2263),
            .I(N__2257));
    InMux I__473 (
            .O(N__2262),
            .I(N__2250));
    InMux I__472 (
            .O(N__2261),
            .I(N__2250));
    InMux I__471 (
            .O(N__2260),
            .I(N__2250));
    Odrv12 I__470 (
            .O(N__2257),
            .I(shift2_0Z0Z_2));
    LocalMux I__469 (
            .O(N__2250),
            .I(shift2_0Z0Z_2));
    CascadeMux I__468 (
            .O(N__2245),
            .I(N__2241));
    InMux I__467 (
            .O(N__2244),
            .I(N__2238));
    InMux I__466 (
            .O(N__2241),
            .I(N__2235));
    LocalMux I__465 (
            .O(N__2238),
            .I(clk_divZ0Z_8));
    LocalMux I__464 (
            .O(N__2235),
            .I(clk_divZ0Z_8));
    InMux I__463 (
            .O(N__2230),
            .I(clk_div_1_cry_7));
    CascadeMux I__462 (
            .O(N__2227),
            .I(N__2223));
    InMux I__461 (
            .O(N__2226),
            .I(N__2220));
    InMux I__460 (
            .O(N__2223),
            .I(N__2217));
    LocalMux I__459 (
            .O(N__2220),
            .I(clk_divZ0Z_9));
    LocalMux I__458 (
            .O(N__2217),
            .I(clk_divZ0Z_9));
    InMux I__457 (
            .O(N__2212),
            .I(bfn_2_9_0_));
    InMux I__456 (
            .O(N__2209),
            .I(clk_div_1_cry_9));
    InMux I__455 (
            .O(N__2206),
            .I(N__2202));
    InMux I__454 (
            .O(N__2205),
            .I(N__2199));
    LocalMux I__453 (
            .O(N__2202),
            .I(clk_divZ0Z_10));
    LocalMux I__452 (
            .O(N__2199),
            .I(clk_divZ0Z_10));
    ClkMux I__451 (
            .O(N__2194),
            .I(N__2161));
    ClkMux I__450 (
            .O(N__2193),
            .I(N__2161));
    ClkMux I__449 (
            .O(N__2192),
            .I(N__2161));
    ClkMux I__448 (
            .O(N__2191),
            .I(N__2161));
    ClkMux I__447 (
            .O(N__2190),
            .I(N__2161));
    ClkMux I__446 (
            .O(N__2189),
            .I(N__2161));
    ClkMux I__445 (
            .O(N__2188),
            .I(N__2161));
    ClkMux I__444 (
            .O(N__2187),
            .I(N__2161));
    ClkMux I__443 (
            .O(N__2186),
            .I(N__2161));
    ClkMux I__442 (
            .O(N__2185),
            .I(N__2161));
    ClkMux I__441 (
            .O(N__2184),
            .I(N__2161));
    GlobalMux I__440 (
            .O(N__2161),
            .I(N__2158));
    gio2CtrlBuf I__439 (
            .O(N__2158),
            .I(CLK_0_c_g));
    InMux I__438 (
            .O(N__2155),
            .I(N__2152));
    LocalMux I__437 (
            .O(N__2152),
            .I(N__2149));
    Span4Mux_s3_h I__436 (
            .O(N__2149),
            .I(N__2145));
    InMux I__435 (
            .O(N__2148),
            .I(N__2142));
    Odrv4 I__434 (
            .O(N__2145),
            .I(upZ0Z_2));
    LocalMux I__433 (
            .O(N__2142),
            .I(upZ0Z_2));
    InMux I__432 (
            .O(N__2137),
            .I(N__2134));
    LocalMux I__431 (
            .O(N__2134),
            .I(N__2130));
    InMux I__430 (
            .O(N__2133),
            .I(N__2127));
    Span4Mux_v I__429 (
            .O(N__2130),
            .I(N__2120));
    LocalMux I__428 (
            .O(N__2127),
            .I(N__2120));
    InMux I__427 (
            .O(N__2126),
            .I(N__2115));
    InMux I__426 (
            .O(N__2125),
            .I(N__2115));
    Odrv4 I__425 (
            .O(N__2120),
            .I(upZ0Z_1));
    LocalMux I__424 (
            .O(N__2115),
            .I(upZ0Z_1));
    CEMux I__423 (
            .O(N__2110),
            .I(N__2107));
    LocalMux I__422 (
            .O(N__2107),
            .I(N__2104));
    Span4Mux_v I__421 (
            .O(N__2104),
            .I(N__2101));
    Odrv4 I__420 (
            .O(N__2101),
            .I(shift_ret_1_RNI69IQZ0));
    InMux I__419 (
            .O(N__2098),
            .I(N__2092));
    InMux I__418 (
            .O(N__2097),
            .I(N__2087));
    InMux I__417 (
            .O(N__2096),
            .I(N__2087));
    InMux I__416 (
            .O(N__2095),
            .I(N__2084));
    LocalMux I__415 (
            .O(N__2092),
            .I(N__2079));
    LocalMux I__414 (
            .O(N__2087),
            .I(N__2079));
    LocalMux I__413 (
            .O(N__2084),
            .I(clk_div_RNI06L91Z0Z_11));
    Odrv4 I__412 (
            .O(N__2079),
            .I(clk_div_RNI06L91Z0Z_11));
    InMux I__411 (
            .O(N__2074),
            .I(N__2068));
    InMux I__410 (
            .O(N__2073),
            .I(N__2063));
    InMux I__409 (
            .O(N__2072),
            .I(N__2063));
    InMux I__408 (
            .O(N__2071),
            .I(N__2060));
    LocalMux I__407 (
            .O(N__2068),
            .I(clk_div_i_11));
    LocalMux I__406 (
            .O(N__2063),
            .I(clk_div_i_11));
    LocalMux I__405 (
            .O(N__2060),
            .I(clk_div_i_11));
    InMux I__404 (
            .O(N__2053),
            .I(N__2048));
    InMux I__403 (
            .O(N__2052),
            .I(N__2045));
    InMux I__402 (
            .O(N__2051),
            .I(N__2042));
    LocalMux I__401 (
            .O(N__2048),
            .I(clk_divZ0Z_1));
    LocalMux I__400 (
            .O(N__2045),
            .I(clk_divZ0Z_1));
    LocalMux I__399 (
            .O(N__2042),
            .I(clk_divZ0Z_1));
    CascadeMux I__398 (
            .O(N__2035),
            .I(N__2029));
    CascadeMux I__397 (
            .O(N__2034),
            .I(N__2026));
    InMux I__396 (
            .O(N__2033),
            .I(N__2023));
    InMux I__395 (
            .O(N__2032),
            .I(N__2020));
    InMux I__394 (
            .O(N__2029),
            .I(N__2017));
    InMux I__393 (
            .O(N__2026),
            .I(N__2014));
    LocalMux I__392 (
            .O(N__2023),
            .I(clk_divZ0Z_0));
    LocalMux I__391 (
            .O(N__2020),
            .I(clk_divZ0Z_0));
    LocalMux I__390 (
            .O(N__2017),
            .I(clk_divZ0Z_0));
    LocalMux I__389 (
            .O(N__2014),
            .I(clk_divZ0Z_0));
    CascadeMux I__388 (
            .O(N__2005),
            .I(N__2001));
    InMux I__387 (
            .O(N__2004),
            .I(N__1998));
    InMux I__386 (
            .O(N__2001),
            .I(N__1995));
    LocalMux I__385 (
            .O(N__1998),
            .I(clk_divZ0Z_2));
    LocalMux I__384 (
            .O(N__1995),
            .I(clk_divZ0Z_2));
    InMux I__383 (
            .O(N__1990),
            .I(clk_div_1_cry_1));
    CascadeMux I__382 (
            .O(N__1987),
            .I(N__1983));
    InMux I__381 (
            .O(N__1986),
            .I(N__1980));
    InMux I__380 (
            .O(N__1983),
            .I(N__1977));
    LocalMux I__379 (
            .O(N__1980),
            .I(clk_divZ0Z_3));
    LocalMux I__378 (
            .O(N__1977),
            .I(clk_divZ0Z_3));
    InMux I__377 (
            .O(N__1972),
            .I(clk_div_1_cry_2));
    CascadeMux I__376 (
            .O(N__1969),
            .I(N__1965));
    InMux I__375 (
            .O(N__1968),
            .I(N__1962));
    InMux I__374 (
            .O(N__1965),
            .I(N__1959));
    LocalMux I__373 (
            .O(N__1962),
            .I(clk_divZ0Z_4));
    LocalMux I__372 (
            .O(N__1959),
            .I(clk_divZ0Z_4));
    InMux I__371 (
            .O(N__1954),
            .I(clk_div_1_cry_3));
    CascadeMux I__370 (
            .O(N__1951),
            .I(N__1947));
    InMux I__369 (
            .O(N__1950),
            .I(N__1944));
    InMux I__368 (
            .O(N__1947),
            .I(N__1941));
    LocalMux I__367 (
            .O(N__1944),
            .I(clk_divZ0Z_5));
    LocalMux I__366 (
            .O(N__1941),
            .I(clk_divZ0Z_5));
    InMux I__365 (
            .O(N__1936),
            .I(clk_div_1_cry_4));
    CascadeMux I__364 (
            .O(N__1933),
            .I(N__1929));
    InMux I__363 (
            .O(N__1932),
            .I(N__1926));
    InMux I__362 (
            .O(N__1929),
            .I(N__1923));
    LocalMux I__361 (
            .O(N__1926),
            .I(clk_divZ0Z_6));
    LocalMux I__360 (
            .O(N__1923),
            .I(clk_divZ0Z_6));
    InMux I__359 (
            .O(N__1918),
            .I(clk_div_1_cry_5));
    CascadeMux I__358 (
            .O(N__1915),
            .I(N__1911));
    InMux I__357 (
            .O(N__1914),
            .I(N__1908));
    InMux I__356 (
            .O(N__1911),
            .I(N__1905));
    LocalMux I__355 (
            .O(N__1908),
            .I(clk_divZ0Z_7));
    LocalMux I__354 (
            .O(N__1905),
            .I(clk_divZ0Z_7));
    InMux I__353 (
            .O(N__1900),
            .I(clk_div_1_cry_6));
    SRMux I__352 (
            .O(N__1897),
            .I(N__1894));
    LocalMux I__351 (
            .O(N__1894),
            .I(N__1890));
    SRMux I__350 (
            .O(N__1893),
            .I(N__1887));
    Span4Mux_s1_h I__349 (
            .O(N__1890),
            .I(N__1882));
    LocalMux I__348 (
            .O(N__1887),
            .I(N__1882));
    Odrv4 I__347 (
            .O(N__1882),
            .I(PWM_NUM_RNIKTNT2Z0Z_0));
    CascadeMux I__346 (
            .O(N__1879),
            .I(PWM_NUM_RNIKTNT2Z0Z_0_cascade_));
    CEMux I__345 (
            .O(N__1876),
            .I(N__1873));
    LocalMux I__344 (
            .O(N__1873),
            .I(N_78_0));
    InMux I__343 (
            .O(N__1870),
            .I(N__1866));
    InMux I__342 (
            .O(N__1869),
            .I(N__1863));
    LocalMux I__341 (
            .O(N__1866),
            .I(PWM_NUMZ0Z_4));
    LocalMux I__340 (
            .O(N__1863),
            .I(PWM_NUMZ0Z_4));
    InMux I__339 (
            .O(N__1858),
            .I(N__1855));
    LocalMux I__338 (
            .O(N__1855),
            .I(g0_3));
    CascadeMux I__337 (
            .O(N__1852),
            .I(N__1846));
    CascadeMux I__336 (
            .O(N__1851),
            .I(N__1843));
    CascadeMux I__335 (
            .O(N__1850),
            .I(N__1840));
    CascadeMux I__334 (
            .O(N__1849),
            .I(N__1837));
    InMux I__333 (
            .O(N__1846),
            .I(N__1833));
    InMux I__332 (
            .O(N__1843),
            .I(N__1828));
    InMux I__331 (
            .O(N__1840),
            .I(N__1828));
    InMux I__330 (
            .O(N__1837),
            .I(N__1825));
    InMux I__329 (
            .O(N__1836),
            .I(N__1822));
    LocalMux I__328 (
            .O(N__1833),
            .I(cntrZ0Z_4));
    LocalMux I__327 (
            .O(N__1828),
            .I(cntrZ0Z_4));
    LocalMux I__326 (
            .O(N__1825),
            .I(cntrZ0Z_4));
    LocalMux I__325 (
            .O(N__1822),
            .I(cntrZ0Z_4));
    CEMux I__324 (
            .O(N__1813),
            .I(N__1810));
    LocalMux I__323 (
            .O(N__1810),
            .I(N__1805));
    CEMux I__322 (
            .O(N__1809),
            .I(N__1802));
    CEMux I__321 (
            .O(N__1808),
            .I(N__1799));
    Span4Mux_v I__320 (
            .O(N__1805),
            .I(N__1794));
    LocalMux I__319 (
            .O(N__1802),
            .I(N__1794));
    LocalMux I__318 (
            .O(N__1799),
            .I(N__1786));
    Span4Mux_h I__317 (
            .O(N__1794),
            .I(N__1783));
    InMux I__316 (
            .O(N__1793),
            .I(N__1774));
    InMux I__315 (
            .O(N__1792),
            .I(N__1774));
    InMux I__314 (
            .O(N__1791),
            .I(N__1774));
    InMux I__313 (
            .O(N__1790),
            .I(N__1774));
    InMux I__312 (
            .O(N__1789),
            .I(N__1771));
    Odrv4 I__311 (
            .O(N__1786),
            .I(clk_div_RNIM1KP1Z0Z_11));
    Odrv4 I__310 (
            .O(N__1783),
            .I(clk_div_RNIM1KP1Z0Z_11));
    LocalMux I__309 (
            .O(N__1774),
            .I(clk_div_RNIM1KP1Z0Z_11));
    LocalMux I__308 (
            .O(N__1771),
            .I(clk_div_RNIM1KP1Z0Z_11));
    InMux I__307 (
            .O(N__1762),
            .I(N__1758));
    InMux I__306 (
            .O(N__1761),
            .I(N__1753));
    LocalMux I__305 (
            .O(N__1758),
            .I(N__1750));
    InMux I__304 (
            .O(N__1757),
            .I(N__1745));
    InMux I__303 (
            .O(N__1756),
            .I(N__1745));
    LocalMux I__302 (
            .O(N__1753),
            .I(cntrZ0Z_3));
    Odrv4 I__301 (
            .O(N__1750),
            .I(cntrZ0Z_3));
    LocalMux I__300 (
            .O(N__1745),
            .I(cntrZ0Z_3));
    InMux I__299 (
            .O(N__1738),
            .I(N__1732));
    InMux I__298 (
            .O(N__1737),
            .I(N__1729));
    InMux I__297 (
            .O(N__1736),
            .I(N__1726));
    InMux I__296 (
            .O(N__1735),
            .I(N__1723));
    LocalMux I__295 (
            .O(N__1732),
            .I(cntrZ0Z_2));
    LocalMux I__294 (
            .O(N__1729),
            .I(cntrZ0Z_2));
    LocalMux I__293 (
            .O(N__1726),
            .I(cntrZ0Z_2));
    LocalMux I__292 (
            .O(N__1723),
            .I(cntrZ0Z_2));
    InMux I__291 (
            .O(N__1714),
            .I(N__1707));
    InMux I__290 (
            .O(N__1713),
            .I(N__1702));
    InMux I__289 (
            .O(N__1712),
            .I(N__1702));
    InMux I__288 (
            .O(N__1711),
            .I(N__1699));
    InMux I__287 (
            .O(N__1710),
            .I(N__1696));
    LocalMux I__286 (
            .O(N__1707),
            .I(cntrZ0Z_1));
    LocalMux I__285 (
            .O(N__1702),
            .I(cntrZ0Z_1));
    LocalMux I__284 (
            .O(N__1699),
            .I(cntrZ0Z_1));
    LocalMux I__283 (
            .O(N__1696),
            .I(cntrZ0Z_1));
    InMux I__282 (
            .O(N__1687),
            .I(N__1682));
    InMux I__281 (
            .O(N__1686),
            .I(N__1677));
    InMux I__280 (
            .O(N__1685),
            .I(N__1677));
    LocalMux I__279 (
            .O(N__1682),
            .I(un2_cntr_c4));
    LocalMux I__278 (
            .O(N__1677),
            .I(un2_cntr_c4));
    CascadeMux I__277 (
            .O(N__1672),
            .I(N__1665));
    CascadeMux I__276 (
            .O(N__1671),
            .I(N__1662));
    CascadeMux I__275 (
            .O(N__1670),
            .I(N__1657));
    CascadeMux I__274 (
            .O(N__1669),
            .I(N__1654));
    InMux I__273 (
            .O(N__1668),
            .I(N__1651));
    InMux I__272 (
            .O(N__1665),
            .I(N__1648));
    InMux I__271 (
            .O(N__1662),
            .I(N__1643));
    InMux I__270 (
            .O(N__1661),
            .I(N__1643));
    InMux I__269 (
            .O(N__1660),
            .I(N__1638));
    InMux I__268 (
            .O(N__1657),
            .I(N__1638));
    InMux I__267 (
            .O(N__1654),
            .I(N__1635));
    LocalMux I__266 (
            .O(N__1651),
            .I(cntrZ0Z_0));
    LocalMux I__265 (
            .O(N__1648),
            .I(cntrZ0Z_0));
    LocalMux I__264 (
            .O(N__1643),
            .I(cntrZ0Z_0));
    LocalMux I__263 (
            .O(N__1638),
            .I(cntrZ0Z_0));
    LocalMux I__262 (
            .O(N__1635),
            .I(cntrZ0Z_0));
    InMux I__261 (
            .O(N__1624),
            .I(N__1620));
    InMux I__260 (
            .O(N__1623),
            .I(N__1617));
    LocalMux I__259 (
            .O(N__1620),
            .I(N__1612));
    LocalMux I__258 (
            .O(N__1617),
            .I(N__1612));
    Odrv4 I__257 (
            .O(N__1612),
            .I(PWM_NUMZ0Z_0));
    InMux I__256 (
            .O(N__1609),
            .I(N__1606));
    LocalMux I__255 (
            .O(N__1606),
            .I(un1_cntr_0));
    CascadeMux I__254 (
            .O(N__1603),
            .I(N__1597));
    InMux I__253 (
            .O(N__1602),
            .I(N__1594));
    InMux I__252 (
            .O(N__1601),
            .I(N__1591));
    InMux I__251 (
            .O(N__1600),
            .I(N__1588));
    InMux I__250 (
            .O(N__1597),
            .I(N__1585));
    LocalMux I__249 (
            .O(N__1594),
            .I(cntrZ0Z_5));
    LocalMux I__248 (
            .O(N__1591),
            .I(cntrZ0Z_5));
    LocalMux I__247 (
            .O(N__1588),
            .I(cntrZ0Z_5));
    LocalMux I__246 (
            .O(N__1585),
            .I(cntrZ0Z_5));
    InMux I__245 (
            .O(N__1576),
            .I(N__1573));
    LocalMux I__244 (
            .O(N__1573),
            .I(N__1569));
    InMux I__243 (
            .O(N__1572),
            .I(N__1566));
    Odrv4 I__242 (
            .O(N__1569),
            .I(PWM_NUMZ0Z_5));
    LocalMux I__241 (
            .O(N__1566),
            .I(PWM_NUMZ0Z_5));
    CascadeMux I__240 (
            .O(N__1561),
            .I(N__1557));
    CascadeMux I__239 (
            .O(N__1560),
            .I(N__1553));
    InMux I__238 (
            .O(N__1557),
            .I(N__1550));
    InMux I__237 (
            .O(N__1556),
            .I(N__1545));
    InMux I__236 (
            .O(N__1553),
            .I(N__1545));
    LocalMux I__235 (
            .O(N__1550),
            .I(cntrZ0Z_6));
    LocalMux I__234 (
            .O(N__1545),
            .I(cntrZ0Z_6));
    IoInMux I__233 (
            .O(N__1540),
            .I(N__1537));
    LocalMux I__232 (
            .O(N__1537),
            .I(N__1534));
    Span12Mux_s1_h I__231 (
            .O(N__1534),
            .I(N__1529));
    InMux I__230 (
            .O(N__1533),
            .I(N__1526));
    InMux I__229 (
            .O(N__1532),
            .I(N__1523));
    Odrv12 I__228 (
            .O(N__1529),
            .I(PORT1_c));
    LocalMux I__227 (
            .O(N__1526),
            .I(PORT1_c));
    LocalMux I__226 (
            .O(N__1523),
            .I(PORT1_c));
    CascadeMux I__225 (
            .O(N__1516),
            .I(N__1513));
    InMux I__224 (
            .O(N__1513),
            .I(N__1510));
    LocalMux I__223 (
            .O(N__1510),
            .I(N__1507));
    Odrv4 I__222 (
            .O(N__1507),
            .I(PORT_r3_1));
    InMux I__221 (
            .O(N__1504),
            .I(N__1498));
    InMux I__220 (
            .O(N__1503),
            .I(N__1498));
    LocalMux I__219 (
            .O(N__1498),
            .I(PWM_NUMZ0Z_3));
    CascadeMux I__218 (
            .O(N__1495),
            .I(N__1492));
    InMux I__217 (
            .O(N__1492),
            .I(N__1489));
    LocalMux I__216 (
            .O(N__1489),
            .I(PWM_NUMZ0Z_1));
    InMux I__215 (
            .O(N__1486),
            .I(N__1473));
    InMux I__214 (
            .O(N__1485),
            .I(N__1473));
    InMux I__213 (
            .O(N__1484),
            .I(N__1473));
    InMux I__212 (
            .O(N__1483),
            .I(N__1473));
    InMux I__211 (
            .O(N__1482),
            .I(N__1470));
    LocalMux I__210 (
            .O(N__1473),
            .I(howZ0Z_0));
    LocalMux I__209 (
            .O(N__1470),
            .I(howZ0Z_0));
    InMux I__208 (
            .O(N__1465),
            .I(N__1449));
    InMux I__207 (
            .O(N__1464),
            .I(N__1449));
    InMux I__206 (
            .O(N__1463),
            .I(N__1449));
    InMux I__205 (
            .O(N__1462),
            .I(N__1449));
    InMux I__204 (
            .O(N__1461),
            .I(N__1449));
    InMux I__203 (
            .O(N__1460),
            .I(N__1446));
    LocalMux I__202 (
            .O(N__1449),
            .I(howZ0Z_2));
    LocalMux I__201 (
            .O(N__1446),
            .I(howZ0Z_2));
    InMux I__200 (
            .O(N__1441),
            .I(N__1428));
    InMux I__199 (
            .O(N__1440),
            .I(N__1428));
    InMux I__198 (
            .O(N__1439),
            .I(N__1428));
    InMux I__197 (
            .O(N__1438),
            .I(N__1428));
    InMux I__196 (
            .O(N__1437),
            .I(N__1425));
    LocalMux I__195 (
            .O(N__1428),
            .I(howZ0Z_1));
    LocalMux I__194 (
            .O(N__1425),
            .I(howZ0Z_1));
    InMux I__193 (
            .O(N__1420),
            .I(N__1417));
    LocalMux I__192 (
            .O(N__1417),
            .I(PWM_NUMZ0Z_2));
    InMux I__191 (
            .O(N__1414),
            .I(N__1411));
    LocalMux I__190 (
            .O(N__1411),
            .I(PORT_r3_2));
    InMux I__189 (
            .O(N__1408),
            .I(N__1402));
    InMux I__188 (
            .O(N__1407),
            .I(N__1402));
    LocalMux I__187 (
            .O(N__1402),
            .I(PORT_r3_3));
    InMux I__186 (
            .O(N__1399),
            .I(N__1396));
    LocalMux I__185 (
            .O(N__1396),
            .I(g0_2));
    CascadeMux I__184 (
            .O(N__1393),
            .I(g0_4_cascade_));
    InMux I__183 (
            .O(N__1390),
            .I(N__1386));
    InMux I__182 (
            .O(N__1389),
            .I(N__1383));
    LocalMux I__181 (
            .O(N__1386),
            .I(delayZ0Z_10));
    LocalMux I__180 (
            .O(N__1383),
            .I(delayZ0Z_10));
    CascadeMux I__179 (
            .O(N__1378),
            .I(N__1375));
    InMux I__178 (
            .O(N__1375),
            .I(N__1371));
    InMux I__177 (
            .O(N__1374),
            .I(N__1368));
    LocalMux I__176 (
            .O(N__1371),
            .I(delayZ0Z_8));
    LocalMux I__175 (
            .O(N__1368),
            .I(delayZ0Z_8));
    InMux I__174 (
            .O(N__1363),
            .I(N__1359));
    InMux I__173 (
            .O(N__1362),
            .I(N__1356));
    LocalMux I__172 (
            .O(N__1359),
            .I(delayZ0Z_9));
    LocalMux I__171 (
            .O(N__1356),
            .I(delayZ0Z_9));
    InMux I__170 (
            .O(N__1351),
            .I(N__1347));
    InMux I__169 (
            .O(N__1350),
            .I(N__1344));
    LocalMux I__168 (
            .O(N__1347),
            .I(delayZ0Z_0));
    LocalMux I__167 (
            .O(N__1344),
            .I(delayZ0Z_0));
    InMux I__166 (
            .O(N__1339),
            .I(N__1335));
    InMux I__165 (
            .O(N__1338),
            .I(N__1332));
    LocalMux I__164 (
            .O(N__1335),
            .I(delayZ0Z_3));
    LocalMux I__163 (
            .O(N__1332),
            .I(delayZ0Z_3));
    CascadeMux I__162 (
            .O(N__1327),
            .I(N__1324));
    InMux I__161 (
            .O(N__1324),
            .I(N__1320));
    InMux I__160 (
            .O(N__1323),
            .I(N__1317));
    LocalMux I__159 (
            .O(N__1320),
            .I(delayZ0Z_1));
    LocalMux I__158 (
            .O(N__1317),
            .I(delayZ0Z_1));
    InMux I__157 (
            .O(N__1312),
            .I(N__1308));
    InMux I__156 (
            .O(N__1311),
            .I(N__1305));
    LocalMux I__155 (
            .O(N__1308),
            .I(delayZ0Z_2));
    LocalMux I__154 (
            .O(N__1305),
            .I(delayZ0Z_2));
    InMux I__153 (
            .O(N__1300),
            .I(N__1297));
    LocalMux I__152 (
            .O(N__1297),
            .I(un1_ten_ms_7));
    InMux I__151 (
            .O(N__1294),
            .I(N__1291));
    LocalMux I__150 (
            .O(N__1291),
            .I(un1_ten_ms_9));
    CascadeMux I__149 (
            .O(N__1288),
            .I(un1_ten_ms_8_cascade_));
    InMux I__148 (
            .O(N__1285),
            .I(N__1282));
    LocalMux I__147 (
            .O(N__1282),
            .I(un1_ten_ms_10));
    InMux I__146 (
            .O(N__1279),
            .I(N__1276));
    LocalMux I__145 (
            .O(N__1276),
            .I(how_1_c2));
    InMux I__144 (
            .O(N__1273),
            .I(clk_div_2_cry_10));
    InMux I__143 (
            .O(N__1270),
            .I(N__1266));
    InMux I__142 (
            .O(N__1269),
            .I(N__1263));
    LocalMux I__141 (
            .O(N__1266),
            .I(delayZ0Z_6));
    LocalMux I__140 (
            .O(N__1263),
            .I(delayZ0Z_6));
    InMux I__139 (
            .O(N__1258),
            .I(N__1254));
    InMux I__138 (
            .O(N__1257),
            .I(N__1251));
    LocalMux I__137 (
            .O(N__1254),
            .I(delayZ0Z_5));
    LocalMux I__136 (
            .O(N__1251),
            .I(delayZ0Z_5));
    InMux I__135 (
            .O(N__1246),
            .I(N__1242));
    InMux I__134 (
            .O(N__1245),
            .I(N__1239));
    LocalMux I__133 (
            .O(N__1242),
            .I(delayZ0Z_4));
    LocalMux I__132 (
            .O(N__1239),
            .I(delayZ0Z_4));
    InMux I__131 (
            .O(N__1234),
            .I(N__1230));
    InMux I__130 (
            .O(N__1233),
            .I(N__1227));
    LocalMux I__129 (
            .O(N__1230),
            .I(delayZ0Z_7));
    LocalMux I__128 (
            .O(N__1227),
            .I(delayZ0Z_7));
    InMux I__127 (
            .O(N__1222),
            .I(bfn_1_3_0_));
    InMux I__126 (
            .O(N__1219),
            .I(delay_cry_8));
    InMux I__125 (
            .O(N__1216),
            .I(delay_cry_9));
    InMux I__124 (
            .O(N__1213),
            .I(delay_cry_10));
    InMux I__123 (
            .O(N__1210),
            .I(delay_cry_11));
    InMux I__122 (
            .O(N__1207),
            .I(delay_cry_12));
    InMux I__121 (
            .O(N__1204),
            .I(delay_cry_13));
    InMux I__120 (
            .O(N__1201),
            .I(N__1195));
    InMux I__119 (
            .O(N__1200),
            .I(N__1195));
    LocalMux I__118 (
            .O(N__1195),
            .I(delayZ0Z_14));
    InMux I__117 (
            .O(N__1192),
            .I(N__1186));
    InMux I__116 (
            .O(N__1191),
            .I(N__1186));
    LocalMux I__115 (
            .O(N__1186),
            .I(delayZ0Z_13));
    CascadeMux I__114 (
            .O(N__1183),
            .I(N__1180));
    InMux I__113 (
            .O(N__1180),
            .I(N__1174));
    InMux I__112 (
            .O(N__1179),
            .I(N__1174));
    LocalMux I__111 (
            .O(N__1174),
            .I(delayZ0Z_12));
    InMux I__110 (
            .O(N__1171),
            .I(N__1165));
    InMux I__109 (
            .O(N__1170),
            .I(N__1165));
    LocalMux I__108 (
            .O(N__1165),
            .I(delayZ0Z_11));
    InMux I__107 (
            .O(N__1162),
            .I(bfn_1_2_0_));
    InMux I__106 (
            .O(N__1159),
            .I(delay_cry_0));
    InMux I__105 (
            .O(N__1156),
            .I(delay_cry_1));
    InMux I__104 (
            .O(N__1153),
            .I(delay_cry_2));
    InMux I__103 (
            .O(N__1150),
            .I(delay_cry_3));
    InMux I__102 (
            .O(N__1147),
            .I(delay_cry_4));
    InMux I__101 (
            .O(N__1144),
            .I(delay_cry_5));
    InMux I__100 (
            .O(N__1141),
            .I(delay_cry_6));
    defparam IN_MUX_bfv_1_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_7_0_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(clk_div_2_cry_8),
            .carryinitout(bfn_1_8_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(clk_div_1_cry_8),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_1_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_2_0_));
    defparam IN_MUX_bfv_1_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_3_0_ (
            .carryinitin(delay_cry_7),
            .carryinitout(bfn_1_3_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam delay_0_LC_1_2_0.C_ON=1'b1;
    defparam delay_0_LC_1_2_0.SEQ_MODE=4'b1000;
    defparam delay_0_LC_1_2_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 delay_0_LC_1_2_0 (
            .in0(_gnd_net_),
            .in1(N__1350),
            .in2(_gnd_net_),
            .in3(N__1162),
            .lcout(delayZ0Z_0),
            .ltout(),
            .carryin(bfn_1_2_0_),
            .carryout(delay_cry_0),
            .clk(N__2194),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_1_LC_1_2_1.C_ON=1'b1;
    defparam delay_1_LC_1_2_1.SEQ_MODE=4'b1000;
    defparam delay_1_LC_1_2_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 delay_1_LC_1_2_1 (
            .in0(_gnd_net_),
            .in1(N__1323),
            .in2(_gnd_net_),
            .in3(N__1159),
            .lcout(delayZ0Z_1),
            .ltout(),
            .carryin(delay_cry_0),
            .carryout(delay_cry_1),
            .clk(N__2194),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_2_LC_1_2_2.C_ON=1'b1;
    defparam delay_2_LC_1_2_2.SEQ_MODE=4'b1000;
    defparam delay_2_LC_1_2_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 delay_2_LC_1_2_2 (
            .in0(_gnd_net_),
            .in1(N__1311),
            .in2(_gnd_net_),
            .in3(N__1156),
            .lcout(delayZ0Z_2),
            .ltout(),
            .carryin(delay_cry_1),
            .carryout(delay_cry_2),
            .clk(N__2194),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_3_LC_1_2_3.C_ON=1'b1;
    defparam delay_3_LC_1_2_3.SEQ_MODE=4'b1000;
    defparam delay_3_LC_1_2_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 delay_3_LC_1_2_3 (
            .in0(_gnd_net_),
            .in1(N__1338),
            .in2(_gnd_net_),
            .in3(N__1153),
            .lcout(delayZ0Z_3),
            .ltout(),
            .carryin(delay_cry_2),
            .carryout(delay_cry_3),
            .clk(N__2194),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_4_LC_1_2_4.C_ON=1'b1;
    defparam delay_4_LC_1_2_4.SEQ_MODE=4'b1000;
    defparam delay_4_LC_1_2_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 delay_4_LC_1_2_4 (
            .in0(_gnd_net_),
            .in1(N__1245),
            .in2(_gnd_net_),
            .in3(N__1150),
            .lcout(delayZ0Z_4),
            .ltout(),
            .carryin(delay_cry_3),
            .carryout(delay_cry_4),
            .clk(N__2194),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_5_LC_1_2_5.C_ON=1'b1;
    defparam delay_5_LC_1_2_5.SEQ_MODE=4'b1000;
    defparam delay_5_LC_1_2_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 delay_5_LC_1_2_5 (
            .in0(_gnd_net_),
            .in1(N__1257),
            .in2(_gnd_net_),
            .in3(N__1147),
            .lcout(delayZ0Z_5),
            .ltout(),
            .carryin(delay_cry_4),
            .carryout(delay_cry_5),
            .clk(N__2194),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_6_LC_1_2_6.C_ON=1'b1;
    defparam delay_6_LC_1_2_6.SEQ_MODE=4'b1000;
    defparam delay_6_LC_1_2_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 delay_6_LC_1_2_6 (
            .in0(_gnd_net_),
            .in1(N__1269),
            .in2(_gnd_net_),
            .in3(N__1144),
            .lcout(delayZ0Z_6),
            .ltout(),
            .carryin(delay_cry_5),
            .carryout(delay_cry_6),
            .clk(N__2194),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_7_LC_1_2_7.C_ON=1'b1;
    defparam delay_7_LC_1_2_7.SEQ_MODE=4'b1000;
    defparam delay_7_LC_1_2_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 delay_7_LC_1_2_7 (
            .in0(_gnd_net_),
            .in1(N__1233),
            .in2(_gnd_net_),
            .in3(N__1141),
            .lcout(delayZ0Z_7),
            .ltout(),
            .carryin(delay_cry_6),
            .carryout(delay_cry_7),
            .clk(N__2194),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_8_LC_1_3_0.C_ON=1'b1;
    defparam delay_8_LC_1_3_0.SEQ_MODE=4'b1000;
    defparam delay_8_LC_1_3_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 delay_8_LC_1_3_0 (
            .in0(_gnd_net_),
            .in1(N__1374),
            .in2(_gnd_net_),
            .in3(N__1222),
            .lcout(delayZ0Z_8),
            .ltout(),
            .carryin(bfn_1_3_0_),
            .carryout(delay_cry_8),
            .clk(N__2192),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_9_LC_1_3_1.C_ON=1'b1;
    defparam delay_9_LC_1_3_1.SEQ_MODE=4'b1000;
    defparam delay_9_LC_1_3_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 delay_9_LC_1_3_1 (
            .in0(_gnd_net_),
            .in1(N__1362),
            .in2(_gnd_net_),
            .in3(N__1219),
            .lcout(delayZ0Z_9),
            .ltout(),
            .carryin(delay_cry_8),
            .carryout(delay_cry_9),
            .clk(N__2192),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_10_LC_1_3_2.C_ON=1'b1;
    defparam delay_10_LC_1_3_2.SEQ_MODE=4'b1000;
    defparam delay_10_LC_1_3_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 delay_10_LC_1_3_2 (
            .in0(_gnd_net_),
            .in1(N__1389),
            .in2(_gnd_net_),
            .in3(N__1216),
            .lcout(delayZ0Z_10),
            .ltout(),
            .carryin(delay_cry_9),
            .carryout(delay_cry_10),
            .clk(N__2192),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_11_LC_1_3_3.C_ON=1'b1;
    defparam delay_11_LC_1_3_3.SEQ_MODE=4'b1000;
    defparam delay_11_LC_1_3_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 delay_11_LC_1_3_3 (
            .in0(_gnd_net_),
            .in1(N__1170),
            .in2(_gnd_net_),
            .in3(N__1213),
            .lcout(delayZ0Z_11),
            .ltout(),
            .carryin(delay_cry_10),
            .carryout(delay_cry_11),
            .clk(N__2192),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_12_LC_1_3_4.C_ON=1'b1;
    defparam delay_12_LC_1_3_4.SEQ_MODE=4'b1000;
    defparam delay_12_LC_1_3_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 delay_12_LC_1_3_4 (
            .in0(_gnd_net_),
            .in1(N__1179),
            .in2(_gnd_net_),
            .in3(N__1210),
            .lcout(delayZ0Z_12),
            .ltout(),
            .carryin(delay_cry_11),
            .carryout(delay_cry_12),
            .clk(N__2192),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_13_LC_1_3_5.C_ON=1'b1;
    defparam delay_13_LC_1_3_5.SEQ_MODE=4'b1000;
    defparam delay_13_LC_1_3_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 delay_13_LC_1_3_5 (
            .in0(_gnd_net_),
            .in1(N__1191),
            .in2(_gnd_net_),
            .in3(N__1207),
            .lcout(delayZ0Z_13),
            .ltout(),
            .carryin(delay_cry_12),
            .carryout(delay_cry_13),
            .clk(N__2192),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_14_LC_1_3_6.C_ON=1'b0;
    defparam delay_14_LC_1_3_6.SEQ_MODE=4'b1000;
    defparam delay_14_LC_1_3_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 delay_14_LC_1_3_6 (
            .in0(_gnd_net_),
            .in1(N__1200),
            .in2(_gnd_net_),
            .in3(N__1204),
            .lcout(delayZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2192),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_RNIABQR_14_LC_1_3_7.C_ON=1'b0;
    defparam delay_RNIABQR_14_LC_1_3_7.SEQ_MODE=4'b0000;
    defparam delay_RNIABQR_14_LC_1_3_7.LUT_INIT=16'b0000000000000001;
    LogicCell40 delay_RNIABQR_14_LC_1_3_7 (
            .in0(N__1201),
            .in1(N__1192),
            .in2(N__1183),
            .in3(N__1171),
            .lcout(un1_ten_ms_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_esr_3_LC_1_5_0.C_ON=1'b0;
    defparam cntr_esr_3_LC_1_5_0.SEQ_MODE=4'b1000;
    defparam cntr_esr_3_LC_1_5_0.LUT_INIT=16'b0110101010101010;
    LogicCell40 cntr_esr_3_LC_1_5_0 (
            .in0(N__1761),
            .in1(N__1738),
            .in2(N__1672),
            .in3(N__1714),
            .lcout(cntrZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2189),
            .ce(N__1876),
            .sr(N__1897));
    defparam cntr_2_LC_1_6_0.C_ON=1'b0;
    defparam cntr_2_LC_1_6_0.SEQ_MODE=4'b1000;
    defparam cntr_2_LC_1_6_0.LUT_INIT=16'b0110101010101010;
    LogicCell40 cntr_2_LC_1_6_0 (
            .in0(N__1737),
            .in1(N__1713),
            .in2(N__1671),
            .in3(N__1792),
            .lcout(cntrZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2186),
            .ce(),
            .sr(N__1893));
    defparam cntr_4_LC_1_6_1.C_ON=1'b0;
    defparam cntr_4_LC_1_6_1.SEQ_MODE=4'b1000;
    defparam cntr_4_LC_1_6_1.LUT_INIT=16'b0111100001111000;
    LogicCell40 cntr_4_LC_1_6_1 (
            .in0(N__1791),
            .in1(N__1685),
            .in2(N__1851),
            .in3(_gnd_net_),
            .lcout(cntrZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2186),
            .ce(),
            .sr(N__1893));
    defparam cntr_5_LC_1_6_3.C_ON=1'b0;
    defparam cntr_5_LC_1_6_3.SEQ_MODE=4'b1000;
    defparam cntr_5_LC_1_6_3.LUT_INIT=16'b0110110011001100;
    LogicCell40 cntr_5_LC_1_6_3 (
            .in0(N__1793),
            .in1(N__1601),
            .in2(N__1850),
            .in3(N__1686),
            .lcout(cntrZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2186),
            .ce(),
            .sr(N__1893));
    defparam cntr_1_LC_1_6_4.C_ON=1'b0;
    defparam cntr_1_LC_1_6_4.SEQ_MODE=4'b1000;
    defparam cntr_1_LC_1_6_4.LUT_INIT=16'b0110011011001100;
    LogicCell40 cntr_1_LC_1_6_4 (
            .in0(N__1661),
            .in1(N__1712),
            .in2(_gnd_net_),
            .in3(N__1790),
            .lcout(cntrZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2186),
            .ce(),
            .sr(N__1893));
    defparam cntr_0_LC_1_6_5.C_ON=1'b0;
    defparam cntr_0_LC_1_6_5.SEQ_MODE=4'b1000;
    defparam cntr_0_LC_1_6_5.LUT_INIT=16'b1001100110101010;
    LogicCell40 cntr_0_LC_1_6_5 (
            .in0(N__1668),
            .in1(N__2074),
            .in2(_gnd_net_),
            .in3(N__2098),
            .lcout(cntrZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2186),
            .ce(),
            .sr(N__1893));
    defparam clk_div_RNI91U1_1_LC_1_7_0.C_ON=1'b1;
    defparam clk_div_RNI91U1_1_LC_1_7_0.SEQ_MODE=4'b0000;
    defparam clk_div_RNI91U1_1_LC_1_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNI91U1_1_LC_1_7_0 (
            .in0(_gnd_net_),
            .in1(N__2051),
            .in2(N__2034),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_7_0_),
            .carryout(clk_div_2_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIF3T2_2_LC_1_7_1.C_ON=1'b1;
    defparam clk_div_RNIF3T2_2_LC_1_7_1.SEQ_MODE=4'b0000;
    defparam clk_div_RNIF3T2_2_LC_1_7_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIF3T2_2_LC_1_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2005),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_1),
            .carryout(clk_div_2_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIM6S3_3_LC_1_7_2.C_ON=1'b1;
    defparam clk_div_RNIM6S3_3_LC_1_7_2.SEQ_MODE=4'b0000;
    defparam clk_div_RNIM6S3_3_LC_1_7_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIM6S3_3_LC_1_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1987),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_2),
            .carryout(clk_div_2_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIUAR4_4_LC_1_7_3.C_ON=1'b1;
    defparam clk_div_RNIUAR4_4_LC_1_7_3.SEQ_MODE=4'b0000;
    defparam clk_div_RNIUAR4_4_LC_1_7_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIUAR4_4_LC_1_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1969),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_3),
            .carryout(clk_div_2_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNI7GQ5_5_LC_1_7_4.C_ON=1'b1;
    defparam clk_div_RNI7GQ5_5_LC_1_7_4.SEQ_MODE=4'b0000;
    defparam clk_div_RNI7GQ5_5_LC_1_7_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNI7GQ5_5_LC_1_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1951),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_4),
            .carryout(clk_div_2_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIHMP6_6_LC_1_7_5.C_ON=1'b1;
    defparam clk_div_RNIHMP6_6_LC_1_7_5.SEQ_MODE=4'b0000;
    defparam clk_div_RNIHMP6_6_LC_1_7_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIHMP6_6_LC_1_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1933),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_5),
            .carryout(clk_div_2_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNISTO7_7_LC_1_7_6.C_ON=1'b1;
    defparam clk_div_RNISTO7_7_LC_1_7_6.SEQ_MODE=4'b0000;
    defparam clk_div_RNISTO7_7_LC_1_7_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNISTO7_7_LC_1_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1915),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_6),
            .carryout(clk_div_2_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNI86O8_8_LC_1_7_7.C_ON=1'b1;
    defparam clk_div_RNI86O8_8_LC_1_7_7.SEQ_MODE=4'b0000;
    defparam clk_div_RNI86O8_8_LC_1_7_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNI86O8_8_LC_1_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2245),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_7),
            .carryout(clk_div_2_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNILFN9_9_LC_1_8_0.C_ON=1'b1;
    defparam clk_div_RNILFN9_9_LC_1_8_0.SEQ_MODE=4'b0000;
    defparam clk_div_RNILFN9_9_LC_1_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNILFN9_9_LC_1_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2227),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_8_0_),
            .carryout(clk_div_2_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIAAMP_10_LC_1_8_1.C_ON=1'b1;
    defparam clk_div_RNIAAMP_10_LC_1_8_1.SEQ_MODE=4'b0000;
    defparam clk_div_RNIAAMP_10_LC_1_8_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIAAMP_10_LC_1_8_1 (
            .in0(_gnd_net_),
            .in1(N__2205),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_9),
            .carryout(clk_div_2_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNI06L91_11_LC_1_8_2.C_ON=1'b0;
    defparam clk_div_RNI06L91_11_LC_1_8_2.SEQ_MODE=4'b0000;
    defparam clk_div_RNI06L91_11_LC_1_8_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 clk_div_RNI06L91_11_LC_1_8_2 (
            .in0(_gnd_net_),
            .in1(N__2071),
            .in2(_gnd_net_),
            .in3(N__1273),
            .lcout(clk_div_RNI06L91Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_1_LC_1_8_4.C_ON=1'b0;
    defparam clk_div_1_LC_1_8_4.SEQ_MODE=4'b1000;
    defparam clk_div_1_LC_1_8_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_div_1_LC_1_8_4 (
            .in0(_gnd_net_),
            .in1(N__2033),
            .in2(_gnd_net_),
            .in3(N__2053),
            .lcout(clk_divZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2184),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_RNIKNK01_4_LC_2_2_1.C_ON=1'b0;
    defparam delay_RNIKNK01_4_LC_2_2_1.SEQ_MODE=4'b0000;
    defparam delay_RNIKNK01_4_LC_2_2_1.LUT_INIT=16'b0000000000010001;
    LogicCell40 delay_RNIKNK01_4_LC_2_2_1 (
            .in0(N__1270),
            .in1(N__1258),
            .in2(_gnd_net_),
            .in3(N__1246),
            .lcout(un1_ten_ms_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_RNI5HJ71_10_LC_2_2_2.C_ON=1'b0;
    defparam delay_RNI5HJ71_10_LC_2_2_2.SEQ_MODE=4'b0000;
    defparam delay_RNI5HJ71_10_LC_2_2_2.LUT_INIT=16'b0000000000000001;
    LogicCell40 delay_RNI5HJ71_10_LC_2_2_2 (
            .in0(N__1234),
            .in1(N__1390),
            .in2(N__1378),
            .in3(N__1363),
            .lcout(un1_ten_ms_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_RNI2HGB1_0_LC_2_2_5.C_ON=1'b0;
    defparam delay_RNI2HGB1_0_LC_2_2_5.SEQ_MODE=4'b0000;
    defparam delay_RNI2HGB1_0_LC_2_2_5.LUT_INIT=16'b0000000000000001;
    LogicCell40 delay_RNI2HGB1_0_LC_2_2_5 (
            .in0(N__1351),
            .in1(N__1339),
            .in2(N__1327),
            .in3(N__1312),
            .lcout(),
            .ltout(un1_ten_ms_8_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam delay_RNI55JF4_10_LC_2_2_6.C_ON=1'b0;
    defparam delay_RNI55JF4_10_LC_2_2_6.SEQ_MODE=4'b0000;
    defparam delay_RNI55JF4_10_LC_2_2_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 delay_RNI55JF4_10_LC_2_2_6 (
            .in0(N__1300),
            .in1(N__1294),
            .in2(N__1288),
            .in3(N__1285),
            .lcout(un1_ten_ms_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam how_RNO_0_2_LC_2_3_6.C_ON=1'b0;
    defparam how_RNO_0_2_LC_2_3_6.SEQ_MODE=4'b0000;
    defparam how_RNO_0_2_LC_2_3_6.LUT_INIT=16'b1011001010111011;
    LogicCell40 how_RNO_0_2_LC_2_3_6 (
            .in0(N__2133),
            .in1(N__2499),
            .in2(N__2560),
            .in3(N__2370),
            .lcout(how_1_c2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam how_1_LC_2_4_1.C_ON=1'b0;
    defparam how_1_LC_2_4_1.SEQ_MODE=4'b1000;
    defparam how_1_LC_2_4_1.LUT_INIT=16'b0110001110011100;
    LogicCell40 how_1_LC_2_4_1 (
            .in0(N__2559),
            .in1(N__2137),
            .in2(N__2380),
            .in3(N__2503),
            .lcout(howZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2193),
            .ce(N__1808),
            .sr(_gnd_net_));
    defparam how_0_LC_2_4_2.C_ON=1'b0;
    defparam how_0_LC_2_4_2.SEQ_MODE=4'b1000;
    defparam how_0_LC_2_4_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 how_0_LC_2_4_2 (
            .in0(_gnd_net_),
            .in1(N__2558),
            .in2(_gnd_net_),
            .in3(N__2376),
            .lcout(howZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2193),
            .ce(N__1808),
            .sr(_gnd_net_));
    defparam PWM_NUM_0_LC_2_4_3.C_ON=1'b0;
    defparam PWM_NUM_0_LC_2_4_3.SEQ_MODE=4'b1000;
    defparam PWM_NUM_0_LC_2_4_3.LUT_INIT=16'b1100110000110011;
    LogicCell40 PWM_NUM_0_LC_2_4_3 (
            .in0(_gnd_net_),
            .in1(N__1460),
            .in2(_gnd_net_),
            .in3(N__1482),
            .lcout(PWM_NUMZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2193),
            .ce(N__1808),
            .sr(_gnd_net_));
    defparam how_2_LC_2_4_4.C_ON=1'b0;
    defparam how_2_LC_2_4_4.SEQ_MODE=4'b1000;
    defparam how_2_LC_2_4_4.LUT_INIT=16'b0110011010011001;
    LogicCell40 how_2_LC_2_4_4 (
            .in0(N__1279),
            .in1(N__2155),
            .in2(_gnd_net_),
            .in3(N__2473),
            .lcout(howZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2193),
            .ce(N__1808),
            .sr(_gnd_net_));
    defparam PORT_r_RNO_1_LC_2_5_0.C_ON=1'b0;
    defparam PORT_r_RNO_1_LC_2_5_0.SEQ_MODE=4'b0000;
    defparam PORT_r_RNO_1_LC_2_5_0.LUT_INIT=16'b1000001001000001;
    LogicCell40 PORT_r_RNO_1_LC_2_5_0 (
            .in0(N__1757),
            .in1(N__1870),
            .in2(N__1849),
            .in3(N__1504),
            .lcout(PORT_r3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam PWM_NUM_3_LC_2_5_1.C_ON=1'b0;
    defparam PWM_NUM_3_LC_2_5_1.SEQ_MODE=4'b1000;
    defparam PWM_NUM_3_LC_2_5_1.LUT_INIT=16'b0000000010001000;
    LogicCell40 PWM_NUM_3_LC_2_5_1 (
            .in0(N__1485),
            .in1(N__1464),
            .in2(_gnd_net_),
            .in3(N__1440),
            .lcout(PWM_NUMZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2191),
            .ce(N__1813),
            .sr(_gnd_net_));
    defparam PWM_NUM_RNIDRQK_3_LC_2_5_2.C_ON=1'b0;
    defparam PWM_NUM_RNIDRQK_3_LC_2_5_2.SEQ_MODE=4'b0000;
    defparam PWM_NUM_RNIDRQK_3_LC_2_5_2.LUT_INIT=16'b1000001001000001;
    LogicCell40 PWM_NUM_RNIDRQK_3_LC_2_5_2 (
            .in0(N__1756),
            .in1(N__1572),
            .in2(N__1603),
            .in3(N__1503),
            .lcout(g0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam PWM_NUM_5_LC_2_5_3.C_ON=1'b0;
    defparam PWM_NUM_5_LC_2_5_3.SEQ_MODE=4'b1000;
    defparam PWM_NUM_5_LC_2_5_3.LUT_INIT=16'b1000100000000000;
    LogicCell40 PWM_NUM_5_LC_2_5_3 (
            .in0(N__1486),
            .in1(N__1465),
            .in2(_gnd_net_),
            .in3(N__1441),
            .lcout(PWM_NUMZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2191),
            .ce(N__1813),
            .sr(_gnd_net_));
    defparam PWM_NUM_4_LC_2_5_4.C_ON=1'b0;
    defparam PWM_NUM_4_LC_2_5_4.SEQ_MODE=4'b1000;
    defparam PWM_NUM_4_LC_2_5_4.LUT_INIT=16'b1000100010001000;
    LogicCell40 PWM_NUM_4_LC_2_5_4 (
            .in0(N__1461),
            .in1(N__1437),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PWM_NUMZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2191),
            .ce(N__1813),
            .sr(_gnd_net_));
    defparam PWM_NUM_1_LC_2_5_5.C_ON=1'b0;
    defparam PWM_NUM_1_LC_2_5_5.SEQ_MODE=4'b1000;
    defparam PWM_NUM_1_LC_2_5_5.LUT_INIT=16'b0001000101100110;
    LogicCell40 PWM_NUM_1_LC_2_5_5 (
            .in0(N__1483),
            .in1(N__1462),
            .in2(_gnd_net_),
            .in3(N__1438),
            .lcout(PWM_NUMZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2191),
            .ce(N__1813),
            .sr(_gnd_net_));
    defparam PWM_NUM_RNIQIR6_1_LC_2_5_6.C_ON=1'b0;
    defparam PWM_NUM_RNIQIR6_1_LC_2_5_6.SEQ_MODE=4'b0000;
    defparam PWM_NUM_RNIQIR6_1_LC_2_5_6.LUT_INIT=16'b1000001001000001;
    LogicCell40 PWM_NUM_RNIQIR6_1_LC_2_5_6 (
            .in0(N__1735),
            .in1(N__1710),
            .in2(N__1495),
            .in3(N__1420),
            .lcout(PORT_r3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam PWM_NUM_2_LC_2_5_7.C_ON=1'b0;
    defparam PWM_NUM_2_LC_2_5_7.SEQ_MODE=4'b1000;
    defparam PWM_NUM_2_LC_2_5_7.LUT_INIT=16'b0110011001000100;
    LogicCell40 PWM_NUM_2_LC_2_5_7 (
            .in0(N__1484),
            .in1(N__1463),
            .in2(_gnd_net_),
            .in3(N__1439),
            .lcout(PWM_NUMZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2191),
            .ce(N__1813),
            .sr(_gnd_net_));
    defparam PORT_r_LC_2_6_0.C_ON=1'b0;
    defparam PORT_r_LC_2_6_0.SEQ_MODE=4'b1000;
    defparam PORT_r_LC_2_6_0.LUT_INIT=16'b0000000010000000;
    LogicCell40 PORT_r_LC_2_6_0 (
            .in0(N__1408),
            .in1(N__1414),
            .in2(N__1516),
            .in3(N__1609),
            .lcout(PORT1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2190),
            .ce(N__1809),
            .sr(_gnd_net_));
    defparam PWM_NUM_RNIQ48Q_0_LC_2_6_1.C_ON=1'b0;
    defparam PWM_NUM_RNIQ48Q_0_LC_2_6_1.SEQ_MODE=4'b0000;
    defparam PWM_NUM_RNIQ48Q_0_LC_2_6_1.LUT_INIT=16'b0010000100000000;
    LogicCell40 PWM_NUM_RNIQ48Q_0_LC_2_6_1 (
            .in0(N__1623),
            .in1(N__2072),
            .in2(N__1669),
            .in3(N__1407),
            .lcout(),
            .ltout(g0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam PWM_NUM_RNIKTNT2_0_LC_2_6_2.C_ON=1'b0;
    defparam PWM_NUM_RNIKTNT2_0_LC_2_6_2.SEQ_MODE=4'b0000;
    defparam PWM_NUM_RNIKTNT2_0_LC_2_6_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 PWM_NUM_RNIKTNT2_0_LC_2_6_2 (
            .in0(N__1858),
            .in1(N__1399),
            .in2(N__1393),
            .in3(N__2097),
            .lcout(PWM_NUM_RNIKTNT2Z0Z_0),
            .ltout(PWM_NUM_RNIKTNT2Z0Z_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_esr_RNO_0_3_LC_2_6_3.C_ON=1'b0;
    defparam cntr_esr_RNO_0_3_LC_2_6_3.SEQ_MODE=4'b0000;
    defparam cntr_esr_RNO_0_3_LC_2_6_3.LUT_INIT=16'b1111111111110000;
    LogicCell40 cntr_esr_RNO_0_3_LC_2_6_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1879),
            .in3(N__1789),
            .lcout(N_78_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIM1KP1_11_LC_2_6_4.C_ON=1'b0;
    defparam clk_div_RNIM1KP1_11_LC_2_6_4.SEQ_MODE=4'b0000;
    defparam clk_div_RNIM1KP1_11_LC_2_6_4.LUT_INIT=16'b0101010100000000;
    LogicCell40 clk_div_RNIM1KP1_11_LC_2_6_4 (
            .in0(N__2073),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2096),
            .lcout(clk_div_RNIM1KP1Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam PWM_NUM_RNIDNV4_4_LC_2_6_5.C_ON=1'b0;
    defparam PWM_NUM_RNIDNV4_4_LC_2_6_5.SEQ_MODE=4'b0000;
    defparam PWM_NUM_RNIDNV4_4_LC_2_6_5.LUT_INIT=16'b0000000000001001;
    LogicCell40 PWM_NUM_RNIDNV4_4_LC_2_6_5 (
            .in0(N__1869),
            .in1(N__1836),
            .in2(N__1560),
            .in3(N__1532),
            .lcout(g0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_6_LC_2_6_7.C_ON=1'b0;
    defparam cntr_6_LC_2_6_7.SEQ_MODE=4'b1000;
    defparam cntr_6_LC_2_6_7.LUT_INIT=16'b0110101010101010;
    LogicCell40 cntr_6_LC_2_6_7 (
            .in0(N__1556),
            .in1(N__1687),
            .in2(N__1852),
            .in3(N__1602),
            .lcout(cntrZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2190),
            .ce(N__1809),
            .sr(_gnd_net_));
    defparam cntr_RNIB8QE_2_LC_2_7_0.C_ON=1'b0;
    defparam cntr_RNIB8QE_2_LC_2_7_0.SEQ_MODE=4'b0000;
    defparam cntr_RNIB8QE_2_LC_2_7_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 cntr_RNIB8QE_2_LC_2_7_0 (
            .in0(N__1762),
            .in1(N__1736),
            .in2(N__1670),
            .in3(N__1711),
            .lcout(un2_cntr_c4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_0_LC_2_7_1.C_ON=1'b0;
    defparam clk_div_0_LC_2_7_1.SEQ_MODE=4'b1000;
    defparam clk_div_0_LC_2_7_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 clk_div_0_LC_2_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2032),
            .lcout(clk_divZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2187),
            .ce(),
            .sr(_gnd_net_));
    defparam PORT_r_RNO_2_LC_2_7_3.C_ON=1'b0;
    defparam PORT_r_RNO_2_LC_2_7_3.SEQ_MODE=4'b0000;
    defparam PORT_r_RNO_2_LC_2_7_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 PORT_r_RNO_2_LC_2_7_3 (
            .in0(_gnd_net_),
            .in1(N__1660),
            .in2(_gnd_net_),
            .in3(N__1624),
            .lcout(un1_cntr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam PORT_r_RNO_0_LC_2_7_4.C_ON=1'b0;
    defparam PORT_r_RNO_0_LC_2_7_4.SEQ_MODE=4'b0000;
    defparam PORT_r_RNO_0_LC_2_7_4.LUT_INIT=16'b0000000000001001;
    LogicCell40 PORT_r_RNO_0_LC_2_7_4 (
            .in0(N__1600),
            .in1(N__1576),
            .in2(N__1561),
            .in3(N__1533),
            .lcout(PORT_r3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_11_LC_2_7_7.C_ON=1'b0;
    defparam clk_div_11_LC_2_7_7.SEQ_MODE=4'b1000;
    defparam clk_div_11_LC_2_7_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 clk_div_11_LC_2_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2095),
            .lcout(clk_div_i_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2187),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_1_cry_1_c_LC_2_8_0.C_ON=1'b1;
    defparam clk_div_1_cry_1_c_LC_2_8_0.SEQ_MODE=4'b0000;
    defparam clk_div_1_cry_1_c_LC_2_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_1_cry_1_c_LC_2_8_0 (
            .in0(_gnd_net_),
            .in1(N__2052),
            .in2(N__2035),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(clk_div_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_2_LC_2_8_1.C_ON=1'b1;
    defparam clk_div_2_LC_2_8_1.SEQ_MODE=4'b1000;
    defparam clk_div_2_LC_2_8_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_2_LC_2_8_1 (
            .in0(_gnd_net_),
            .in1(N__2004),
            .in2(_gnd_net_),
            .in3(N__1990),
            .lcout(clk_divZ0Z_2),
            .ltout(),
            .carryin(clk_div_1_cry_1),
            .carryout(clk_div_1_cry_2),
            .clk(N__2185),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_3_LC_2_8_2.C_ON=1'b1;
    defparam clk_div_3_LC_2_8_2.SEQ_MODE=4'b1000;
    defparam clk_div_3_LC_2_8_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_3_LC_2_8_2 (
            .in0(_gnd_net_),
            .in1(N__1986),
            .in2(_gnd_net_),
            .in3(N__1972),
            .lcout(clk_divZ0Z_3),
            .ltout(),
            .carryin(clk_div_1_cry_2),
            .carryout(clk_div_1_cry_3),
            .clk(N__2185),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_4_LC_2_8_3.C_ON=1'b1;
    defparam clk_div_4_LC_2_8_3.SEQ_MODE=4'b1000;
    defparam clk_div_4_LC_2_8_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_4_LC_2_8_3 (
            .in0(_gnd_net_),
            .in1(N__1968),
            .in2(_gnd_net_),
            .in3(N__1954),
            .lcout(clk_divZ0Z_4),
            .ltout(),
            .carryin(clk_div_1_cry_3),
            .carryout(clk_div_1_cry_4),
            .clk(N__2185),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_5_LC_2_8_4.C_ON=1'b1;
    defparam clk_div_5_LC_2_8_4.SEQ_MODE=4'b1000;
    defparam clk_div_5_LC_2_8_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_5_LC_2_8_4 (
            .in0(_gnd_net_),
            .in1(N__1950),
            .in2(_gnd_net_),
            .in3(N__1936),
            .lcout(clk_divZ0Z_5),
            .ltout(),
            .carryin(clk_div_1_cry_4),
            .carryout(clk_div_1_cry_5),
            .clk(N__2185),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_6_LC_2_8_5.C_ON=1'b1;
    defparam clk_div_6_LC_2_8_5.SEQ_MODE=4'b1000;
    defparam clk_div_6_LC_2_8_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_6_LC_2_8_5 (
            .in0(_gnd_net_),
            .in1(N__1932),
            .in2(_gnd_net_),
            .in3(N__1918),
            .lcout(clk_divZ0Z_6),
            .ltout(),
            .carryin(clk_div_1_cry_5),
            .carryout(clk_div_1_cry_6),
            .clk(N__2185),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_7_LC_2_8_6.C_ON=1'b1;
    defparam clk_div_7_LC_2_8_6.SEQ_MODE=4'b1000;
    defparam clk_div_7_LC_2_8_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_7_LC_2_8_6 (
            .in0(_gnd_net_),
            .in1(N__1914),
            .in2(_gnd_net_),
            .in3(N__1900),
            .lcout(clk_divZ0Z_7),
            .ltout(),
            .carryin(clk_div_1_cry_6),
            .carryout(clk_div_1_cry_7),
            .clk(N__2185),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_8_LC_2_8_7.C_ON=1'b1;
    defparam clk_div_8_LC_2_8_7.SEQ_MODE=4'b1000;
    defparam clk_div_8_LC_2_8_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_8_LC_2_8_7 (
            .in0(_gnd_net_),
            .in1(N__2244),
            .in2(_gnd_net_),
            .in3(N__2230),
            .lcout(clk_divZ0Z_8),
            .ltout(),
            .carryin(clk_div_1_cry_7),
            .carryout(clk_div_1_cry_8),
            .clk(N__2185),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_9_LC_2_9_0.C_ON=1'b1;
    defparam clk_div_9_LC_2_9_0.SEQ_MODE=4'b1000;
    defparam clk_div_9_LC_2_9_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_9_LC_2_9_0 (
            .in0(_gnd_net_),
            .in1(N__2226),
            .in2(_gnd_net_),
            .in3(N__2212),
            .lcout(clk_divZ0Z_9),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(clk_div_1_cry_9),
            .clk(N__2188),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_10_LC_2_9_1.C_ON=1'b0;
    defparam clk_div_10_LC_2_9_1.SEQ_MODE=4'b1000;
    defparam clk_div_10_LC_2_9_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 clk_div_10_LC_2_9_1 (
            .in0(_gnd_net_),
            .in1(N__2206),
            .in2(_gnd_net_),
            .in3(N__2209),
            .lcout(clk_divZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2188),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_ret_1_LC_4_2_0.C_ON=1'b0;
    defparam shift_ret_1_LC_4_2_0.SEQ_MODE=4'b1000;
    defparam shift_ret_1_LC_4_2_0.LUT_INIT=16'b1010000000000000;
    LogicCell40 shift_ret_1_LC_4_2_0 (
            .in0(N__2519),
            .in1(_gnd_net_),
            .in2(N__2632),
            .in3(N__2573),
            .lcout(level_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2309),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_0_2_LC_4_2_3.C_ON=1'b0;
    defparam shift_0_2_LC_4_2_3.SEQ_MODE=4'b1000;
    defparam shift_0_2_LC_4_2_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 shift_0_2_LC_4_2_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2627),
            .lcout(shift_0Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2309),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_0_1_LC_4_2_4.C_ON=1'b0;
    defparam shift_0_1_LC_4_2_4.SEQ_MODE=4'b1000;
    defparam shift_0_1_LC_4_2_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift_0_1_LC_4_2_4 (
            .in0(N__2518),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift_0Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2309),
            .ce(),
            .sr(_gnd_net_));
    defparam shift_ret_1_RNI69IQ_LC_4_2_5.C_ON=1'b0;
    defparam shift_ret_1_RNI69IQ_LC_4_2_5.SEQ_MODE=4'b0000;
    defparam shift_ret_1_RNI69IQ_LC_4_2_5.LUT_INIT=16'b0000100000000000;
    LogicCell40 shift_ret_1_RNI69IQ_LC_4_2_5 (
            .in0(N__2574),
            .in1(N__2520),
            .in2(N__2592),
            .in3(N__2631),
            .lcout(shift_ret_1_RNI69IQZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam up_2_LC_4_3_2.C_ON=1'b0;
    defparam up_2_LC_4_3_2.SEQ_MODE=4'b1000;
    defparam up_2_LC_4_3_2.LUT_INIT=16'b0110011011001100;
    LogicCell40 up_2_LC_4_3_2 (
            .in0(N__2541),
            .in1(N__2148),
            .in2(_gnd_net_),
            .in3(N__2126),
            .lcout(upZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2330),
            .ce(N__2110),
            .sr(_gnd_net_));
    defparam up_1_LC_4_3_5.C_ON=1'b0;
    defparam up_1_LC_4_3_5.SEQ_MODE=4'b1000;
    defparam up_1_LC_4_3_5.LUT_INIT=16'b0101010110101010;
    LogicCell40 up_1_LC_4_3_5 (
            .in0(N__2125),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2540),
            .lcout(upZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2330),
            .ce(N__2110),
            .sr(_gnd_net_));
    defparam up_e_0_LC_5_2_7.C_ON=1'b0;
    defparam up_e_0_LC_5_2_7.SEQ_MODE=4'b1000;
    defparam up_e_0_LC_5_2_7.LUT_INIT=16'b1100011011001100;
    LogicCell40 up_e_0_LC_5_2_7 (
            .in0(N__2626),
            .in1(N__2539),
            .in2(N__2593),
            .in3(N__2575),
            .lcout(upZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2325),
            .ce(N__2521),
            .sr(_gnd_net_));
    defparam down_1_LC_5_3_0.C_ON=1'b0;
    defparam down_1_LC_5_3_0.SEQ_MODE=4'b1000;
    defparam down_1_LC_5_3_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 down_1_LC_5_3_0 (
            .in0(_gnd_net_),
            .in1(N__2491),
            .in2(_gnd_net_),
            .in3(N__2361),
            .lcout(downZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2334),
            .ce(N__2455),
            .sr(_gnd_net_));
    defparam down_2_LC_5_3_2.C_ON=1'b0;
    defparam down_2_LC_5_3_2.SEQ_MODE=4'b1000;
    defparam down_2_LC_5_3_2.LUT_INIT=16'b0110011010101010;
    LogicCell40 down_2_LC_5_3_2 (
            .in0(N__2466),
            .in1(N__2492),
            .in2(_gnd_net_),
            .in3(N__2362),
            .lcout(downZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2334),
            .ce(N__2455),
            .sr(_gnd_net_));
    defparam shift2_0_2_LC_6_2_1.C_ON=1'b0;
    defparam shift2_0_2_LC_6_2_1.SEQ_MODE=4'b1000;
    defparam shift2_0_2_LC_6_2_1.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift2_0_2_LC_6_2_1 (
            .in0(N__2401),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift2_0Z0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2326),
            .ce(),
            .sr(_gnd_net_));
    defparam shift2_ret_1_RNITCI51_LC_6_2_4.C_ON=1'b0;
    defparam shift2_ret_1_RNITCI51_LC_6_2_4.SEQ_MODE=4'b0000;
    defparam shift2_ret_1_RNITCI51_LC_6_2_4.LUT_INIT=16'b0100000000000000;
    LogicCell40 shift2_ret_1_RNITCI51_LC_6_2_4 (
            .in0(N__2439),
            .in1(N__2405),
            .in2(N__2428),
            .in3(N__2262),
            .lcout(shift2_ret_1_RNITCIZ0Z51),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam shift2_ret_1_LC_6_2_5.C_ON=1'b0;
    defparam shift2_ret_1_LC_6_2_5.SEQ_MODE=4'b1000;
    defparam shift2_ret_1_LC_6_2_5.LUT_INIT=16'b1010000000000000;
    LogicCell40 shift2_ret_1_LC_6_2_5 (
            .in0(N__2261),
            .in1(_gnd_net_),
            .in2(N__2409),
            .in3(N__2423),
            .lcout(level2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2326),
            .ce(),
            .sr(_gnd_net_));
    defparam shift2_0_1_LC_6_2_7.C_ON=1'b0;
    defparam shift2_0_1_LC_6_2_7.SEQ_MODE=4'b1000;
    defparam shift2_0_1_LC_6_2_7.LUT_INIT=16'b1010101010101010;
    LogicCell40 shift2_0_1_LC_6_2_7 (
            .in0(N__2260),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(shift2_0Z0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2326),
            .ce(),
            .sr(_gnd_net_));
    defparam down_e_0_LC_6_3_4.C_ON=1'b0;
    defparam down_e_0_LC_6_3_4.SEQ_MODE=4'b1000;
    defparam down_e_0_LC_6_3_4.LUT_INIT=16'b1011010011110000;
    LogicCell40 down_e_0_LC_6_3_4 (
            .in0(N__2440),
            .in1(N__2427),
            .in2(N__2369),
            .in3(N__2410),
            .lcout(downZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2335),
            .ce(N__2269),
            .sr(_gnd_net_));
endmodule // top
