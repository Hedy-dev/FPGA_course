-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jul 13 2021 16:01:58

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    PORT1 : out std_logic;
    CLK : in std_logic;
    BUT2 : in std_logic;
    BUT1 : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__2680\ : std_logic;
signal \N__2679\ : std_logic;
signal \N__2678\ : std_logic;
signal \N__2669\ : std_logic;
signal \N__2668\ : std_logic;
signal \N__2667\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2658\ : std_logic;
signal \N__2651\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2631\ : std_logic;
signal \N__2628\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2619\ : std_logic;
signal \N__2616\ : std_logic;
signal \N__2613\ : std_logic;
signal \N__2610\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2589\ : std_logic;
signal \N__2586\ : std_logic;
signal \N__2583\ : std_logic;
signal \N__2580\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2565\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2559\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2550\ : std_logic;
signal \N__2547\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2539\ : std_logic;
signal \N__2536\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2518\ : std_logic;
signal \N__2515\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2480\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2470\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2466\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2449\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2439\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2423\ : std_logic;
signal \N__2420\ : std_logic;
signal \N__2415\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2405\ : std_logic;
signal \N__2402\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2380\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2370\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2361\ : std_logic;
signal \N__2358\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2352\ : std_logic;
signal \N__2347\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2335\ : std_logic;
signal \N__2334\ : std_logic;
signal \N__2331\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2326\ : std_logic;
signal \N__2325\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2316\ : std_logic;
signal \N__2313\ : std_logic;
signal \N__2310\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2298\ : std_logic;
signal \N__2295\ : std_logic;
signal \N__2292\ : std_logic;
signal \N__2289\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2281\ : std_logic;
signal \N__2278\ : std_logic;
signal \N__2269\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2260\ : std_logic;
signal \N__2257\ : std_logic;
signal \N__2250\ : std_logic;
signal \N__2245\ : std_logic;
signal \N__2244\ : std_logic;
signal \N__2241\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2230\ : std_logic;
signal \N__2227\ : std_logic;
signal \N__2226\ : std_logic;
signal \N__2223\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2212\ : std_logic;
signal \N__2209\ : std_logic;
signal \N__2206\ : std_logic;
signal \N__2205\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2194\ : std_logic;
signal \N__2193\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2191\ : std_logic;
signal \N__2190\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2188\ : std_logic;
signal \N__2187\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2185\ : std_logic;
signal \N__2184\ : std_logic;
signal \N__2161\ : std_logic;
signal \N__2158\ : std_logic;
signal \N__2155\ : std_logic;
signal \N__2152\ : std_logic;
signal \N__2149\ : std_logic;
signal \N__2148\ : std_logic;
signal \N__2145\ : std_logic;
signal \N__2142\ : std_logic;
signal \N__2137\ : std_logic;
signal \N__2134\ : std_logic;
signal \N__2133\ : std_logic;
signal \N__2130\ : std_logic;
signal \N__2127\ : std_logic;
signal \N__2126\ : std_logic;
signal \N__2125\ : std_logic;
signal \N__2120\ : std_logic;
signal \N__2115\ : std_logic;
signal \N__2110\ : std_logic;
signal \N__2107\ : std_logic;
signal \N__2104\ : std_logic;
signal \N__2101\ : std_logic;
signal \N__2098\ : std_logic;
signal \N__2097\ : std_logic;
signal \N__2096\ : std_logic;
signal \N__2095\ : std_logic;
signal \N__2092\ : std_logic;
signal \N__2087\ : std_logic;
signal \N__2084\ : std_logic;
signal \N__2079\ : std_logic;
signal \N__2074\ : std_logic;
signal \N__2073\ : std_logic;
signal \N__2072\ : std_logic;
signal \N__2071\ : std_logic;
signal \N__2068\ : std_logic;
signal \N__2063\ : std_logic;
signal \N__2060\ : std_logic;
signal \N__2053\ : std_logic;
signal \N__2052\ : std_logic;
signal \N__2051\ : std_logic;
signal \N__2048\ : std_logic;
signal \N__2045\ : std_logic;
signal \N__2042\ : std_logic;
signal \N__2035\ : std_logic;
signal \N__2034\ : std_logic;
signal \N__2033\ : std_logic;
signal \N__2032\ : std_logic;
signal \N__2029\ : std_logic;
signal \N__2026\ : std_logic;
signal \N__2023\ : std_logic;
signal \N__2020\ : std_logic;
signal \N__2017\ : std_logic;
signal \N__2014\ : std_logic;
signal \N__2005\ : std_logic;
signal \N__2004\ : std_logic;
signal \N__2001\ : std_logic;
signal \N__1998\ : std_logic;
signal \N__1995\ : std_logic;
signal \N__1990\ : std_logic;
signal \N__1987\ : std_logic;
signal \N__1986\ : std_logic;
signal \N__1983\ : std_logic;
signal \N__1980\ : std_logic;
signal \N__1977\ : std_logic;
signal \N__1972\ : std_logic;
signal \N__1969\ : std_logic;
signal \N__1968\ : std_logic;
signal \N__1965\ : std_logic;
signal \N__1962\ : std_logic;
signal \N__1959\ : std_logic;
signal \N__1954\ : std_logic;
signal \N__1951\ : std_logic;
signal \N__1950\ : std_logic;
signal \N__1947\ : std_logic;
signal \N__1944\ : std_logic;
signal \N__1941\ : std_logic;
signal \N__1936\ : std_logic;
signal \N__1933\ : std_logic;
signal \N__1932\ : std_logic;
signal \N__1929\ : std_logic;
signal \N__1926\ : std_logic;
signal \N__1923\ : std_logic;
signal \N__1918\ : std_logic;
signal \N__1915\ : std_logic;
signal \N__1914\ : std_logic;
signal \N__1911\ : std_logic;
signal \N__1908\ : std_logic;
signal \N__1905\ : std_logic;
signal \N__1900\ : std_logic;
signal \N__1897\ : std_logic;
signal \N__1894\ : std_logic;
signal \N__1893\ : std_logic;
signal \N__1890\ : std_logic;
signal \N__1887\ : std_logic;
signal \N__1882\ : std_logic;
signal \N__1879\ : std_logic;
signal \N__1876\ : std_logic;
signal \N__1873\ : std_logic;
signal \N__1870\ : std_logic;
signal \N__1869\ : std_logic;
signal \N__1866\ : std_logic;
signal \N__1863\ : std_logic;
signal \N__1858\ : std_logic;
signal \N__1855\ : std_logic;
signal \N__1852\ : std_logic;
signal \N__1851\ : std_logic;
signal \N__1850\ : std_logic;
signal \N__1849\ : std_logic;
signal \N__1846\ : std_logic;
signal \N__1843\ : std_logic;
signal \N__1840\ : std_logic;
signal \N__1837\ : std_logic;
signal \N__1836\ : std_logic;
signal \N__1833\ : std_logic;
signal \N__1828\ : std_logic;
signal \N__1825\ : std_logic;
signal \N__1822\ : std_logic;
signal \N__1813\ : std_logic;
signal \N__1810\ : std_logic;
signal \N__1809\ : std_logic;
signal \N__1808\ : std_logic;
signal \N__1805\ : std_logic;
signal \N__1802\ : std_logic;
signal \N__1799\ : std_logic;
signal \N__1794\ : std_logic;
signal \N__1793\ : std_logic;
signal \N__1792\ : std_logic;
signal \N__1791\ : std_logic;
signal \N__1790\ : std_logic;
signal \N__1789\ : std_logic;
signal \N__1786\ : std_logic;
signal \N__1783\ : std_logic;
signal \N__1774\ : std_logic;
signal \N__1771\ : std_logic;
signal \N__1762\ : std_logic;
signal \N__1761\ : std_logic;
signal \N__1758\ : std_logic;
signal \N__1757\ : std_logic;
signal \N__1756\ : std_logic;
signal \N__1753\ : std_logic;
signal \N__1750\ : std_logic;
signal \N__1745\ : std_logic;
signal \N__1738\ : std_logic;
signal \N__1737\ : std_logic;
signal \N__1736\ : std_logic;
signal \N__1735\ : std_logic;
signal \N__1732\ : std_logic;
signal \N__1729\ : std_logic;
signal \N__1726\ : std_logic;
signal \N__1723\ : std_logic;
signal \N__1714\ : std_logic;
signal \N__1713\ : std_logic;
signal \N__1712\ : std_logic;
signal \N__1711\ : std_logic;
signal \N__1710\ : std_logic;
signal \N__1707\ : std_logic;
signal \N__1702\ : std_logic;
signal \N__1699\ : std_logic;
signal \N__1696\ : std_logic;
signal \N__1687\ : std_logic;
signal \N__1686\ : std_logic;
signal \N__1685\ : std_logic;
signal \N__1682\ : std_logic;
signal \N__1677\ : std_logic;
signal \N__1672\ : std_logic;
signal \N__1671\ : std_logic;
signal \N__1670\ : std_logic;
signal \N__1669\ : std_logic;
signal \N__1668\ : std_logic;
signal \N__1665\ : std_logic;
signal \N__1662\ : std_logic;
signal \N__1661\ : std_logic;
signal \N__1660\ : std_logic;
signal \N__1657\ : std_logic;
signal \N__1654\ : std_logic;
signal \N__1651\ : std_logic;
signal \N__1648\ : std_logic;
signal \N__1643\ : std_logic;
signal \N__1638\ : std_logic;
signal \N__1635\ : std_logic;
signal \N__1624\ : std_logic;
signal \N__1623\ : std_logic;
signal \N__1620\ : std_logic;
signal \N__1617\ : std_logic;
signal \N__1612\ : std_logic;
signal \N__1609\ : std_logic;
signal \N__1606\ : std_logic;
signal \N__1603\ : std_logic;
signal \N__1602\ : std_logic;
signal \N__1601\ : std_logic;
signal \N__1600\ : std_logic;
signal \N__1597\ : std_logic;
signal \N__1594\ : std_logic;
signal \N__1591\ : std_logic;
signal \N__1588\ : std_logic;
signal \N__1585\ : std_logic;
signal \N__1576\ : std_logic;
signal \N__1573\ : std_logic;
signal \N__1572\ : std_logic;
signal \N__1569\ : std_logic;
signal \N__1566\ : std_logic;
signal \N__1561\ : std_logic;
signal \N__1560\ : std_logic;
signal \N__1557\ : std_logic;
signal \N__1556\ : std_logic;
signal \N__1553\ : std_logic;
signal \N__1550\ : std_logic;
signal \N__1545\ : std_logic;
signal \N__1540\ : std_logic;
signal \N__1537\ : std_logic;
signal \N__1534\ : std_logic;
signal \N__1533\ : std_logic;
signal \N__1532\ : std_logic;
signal \N__1529\ : std_logic;
signal \N__1526\ : std_logic;
signal \N__1523\ : std_logic;
signal \N__1516\ : std_logic;
signal \N__1513\ : std_logic;
signal \N__1510\ : std_logic;
signal \N__1507\ : std_logic;
signal \N__1504\ : std_logic;
signal \N__1503\ : std_logic;
signal \N__1498\ : std_logic;
signal \N__1495\ : std_logic;
signal \N__1492\ : std_logic;
signal \N__1489\ : std_logic;
signal \N__1486\ : std_logic;
signal \N__1485\ : std_logic;
signal \N__1484\ : std_logic;
signal \N__1483\ : std_logic;
signal \N__1482\ : std_logic;
signal \N__1473\ : std_logic;
signal \N__1470\ : std_logic;
signal \N__1465\ : std_logic;
signal \N__1464\ : std_logic;
signal \N__1463\ : std_logic;
signal \N__1462\ : std_logic;
signal \N__1461\ : std_logic;
signal \N__1460\ : std_logic;
signal \N__1449\ : std_logic;
signal \N__1446\ : std_logic;
signal \N__1441\ : std_logic;
signal \N__1440\ : std_logic;
signal \N__1439\ : std_logic;
signal \N__1438\ : std_logic;
signal \N__1437\ : std_logic;
signal \N__1428\ : std_logic;
signal \N__1425\ : std_logic;
signal \N__1420\ : std_logic;
signal \N__1417\ : std_logic;
signal \N__1414\ : std_logic;
signal \N__1411\ : std_logic;
signal \N__1408\ : std_logic;
signal \N__1407\ : std_logic;
signal \N__1402\ : std_logic;
signal \N__1399\ : std_logic;
signal \N__1396\ : std_logic;
signal \N__1393\ : std_logic;
signal \N__1390\ : std_logic;
signal \N__1389\ : std_logic;
signal \N__1386\ : std_logic;
signal \N__1383\ : std_logic;
signal \N__1378\ : std_logic;
signal \N__1375\ : std_logic;
signal \N__1374\ : std_logic;
signal \N__1371\ : std_logic;
signal \N__1368\ : std_logic;
signal \N__1363\ : std_logic;
signal \N__1362\ : std_logic;
signal \N__1359\ : std_logic;
signal \N__1356\ : std_logic;
signal \N__1351\ : std_logic;
signal \N__1350\ : std_logic;
signal \N__1347\ : std_logic;
signal \N__1344\ : std_logic;
signal \N__1339\ : std_logic;
signal \N__1338\ : std_logic;
signal \N__1335\ : std_logic;
signal \N__1332\ : std_logic;
signal \N__1327\ : std_logic;
signal \N__1324\ : std_logic;
signal \N__1323\ : std_logic;
signal \N__1320\ : std_logic;
signal \N__1317\ : std_logic;
signal \N__1312\ : std_logic;
signal \N__1311\ : std_logic;
signal \N__1308\ : std_logic;
signal \N__1305\ : std_logic;
signal \N__1300\ : std_logic;
signal \N__1297\ : std_logic;
signal \N__1294\ : std_logic;
signal \N__1291\ : std_logic;
signal \N__1288\ : std_logic;
signal \N__1285\ : std_logic;
signal \N__1282\ : std_logic;
signal \N__1279\ : std_logic;
signal \N__1276\ : std_logic;
signal \N__1273\ : std_logic;
signal \N__1270\ : std_logic;
signal \N__1269\ : std_logic;
signal \N__1266\ : std_logic;
signal \N__1263\ : std_logic;
signal \N__1258\ : std_logic;
signal \N__1257\ : std_logic;
signal \N__1254\ : std_logic;
signal \N__1251\ : std_logic;
signal \N__1246\ : std_logic;
signal \N__1245\ : std_logic;
signal \N__1242\ : std_logic;
signal \N__1239\ : std_logic;
signal \N__1234\ : std_logic;
signal \N__1233\ : std_logic;
signal \N__1230\ : std_logic;
signal \N__1227\ : std_logic;
signal \N__1222\ : std_logic;
signal \N__1219\ : std_logic;
signal \N__1216\ : std_logic;
signal \N__1213\ : std_logic;
signal \N__1210\ : std_logic;
signal \N__1207\ : std_logic;
signal \N__1204\ : std_logic;
signal \N__1201\ : std_logic;
signal \N__1200\ : std_logic;
signal \N__1195\ : std_logic;
signal \N__1192\ : std_logic;
signal \N__1191\ : std_logic;
signal \N__1186\ : std_logic;
signal \N__1183\ : std_logic;
signal \N__1180\ : std_logic;
signal \N__1179\ : std_logic;
signal \N__1174\ : std_logic;
signal \N__1171\ : std_logic;
signal \N__1170\ : std_logic;
signal \N__1165\ : std_logic;
signal \N__1162\ : std_logic;
signal \N__1159\ : std_logic;
signal \N__1156\ : std_logic;
signal \N__1153\ : std_logic;
signal \N__1150\ : std_logic;
signal \N__1147\ : std_logic;
signal \N__1144\ : std_logic;
signal \N__1141\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_1_2_0_\ : std_logic;
signal delay_cry_0 : std_logic;
signal delay_cry_1 : std_logic;
signal delay_cry_2 : std_logic;
signal delay_cry_3 : std_logic;
signal delay_cry_4 : std_logic;
signal delay_cry_5 : std_logic;
signal delay_cry_6 : std_logic;
signal delay_cry_7 : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal delay_cry_8 : std_logic;
signal delay_cry_9 : std_logic;
signal delay_cry_10 : std_logic;
signal delay_cry_11 : std_logic;
signal delay_cry_12 : std_logic;
signal delay_cry_13 : std_logic;
signal \delayZ0Z_14\ : std_logic;
signal \delayZ0Z_13\ : std_logic;
signal \delayZ0Z_12\ : std_logic;
signal \delayZ0Z_11\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal clk_div_2_cry_1 : std_logic;
signal clk_div_2_cry_2 : std_logic;
signal clk_div_2_cry_3 : std_logic;
signal clk_div_2_cry_4 : std_logic;
signal clk_div_2_cry_5 : std_logic;
signal clk_div_2_cry_6 : std_logic;
signal clk_div_2_cry_7 : std_logic;
signal clk_div_2_cry_8 : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal clk_div_2_cry_9 : std_logic;
signal clk_div_2_cry_10 : std_logic;
signal \delayZ0Z_6\ : std_logic;
signal \delayZ0Z_5\ : std_logic;
signal \delayZ0Z_4\ : std_logic;
signal \delayZ0Z_7\ : std_logic;
signal \delayZ0Z_10\ : std_logic;
signal \delayZ0Z_8\ : std_logic;
signal \delayZ0Z_9\ : std_logic;
signal \delayZ0Z_0\ : std_logic;
signal \delayZ0Z_3\ : std_logic;
signal \delayZ0Z_1\ : std_logic;
signal \delayZ0Z_2\ : std_logic;
signal un1_ten_ms_7 : std_logic;
signal un1_ten_ms_9 : std_logic;
signal \un1_ten_ms_8_cascade_\ : std_logic;
signal un1_ten_ms_10 : std_logic;
signal how_1_c2 : std_logic;
signal \PWM_NUMZ0Z_3\ : std_logic;
signal \PWM_NUMZ0Z_1\ : std_logic;
signal \howZ0Z_0\ : std_logic;
signal \howZ0Z_2\ : std_logic;
signal \howZ0Z_1\ : std_logic;
signal \PWM_NUMZ0Z_2\ : std_logic;
signal \PORT_r3_2\ : std_logic;
signal \PORT_r3_3\ : std_logic;
signal g0_2 : std_logic;
signal \g0_4_cascade_\ : std_logic;
signal \PWM_NUM_RNIKTNT2Z0Z_0\ : std_logic;
signal \PWM_NUM_RNIKTNT2Z0Z_0_cascade_\ : std_logic;
signal \N_78_0\ : std_logic;
signal \PWM_NUMZ0Z_4\ : std_logic;
signal g0_3 : std_logic;
signal \cntrZ0Z_4\ : std_logic;
signal \clk_div_RNIM1KP1Z0Z_11\ : std_logic;
signal \cntrZ0Z_3\ : std_logic;
signal \cntrZ0Z_2\ : std_logic;
signal \cntrZ0Z_1\ : std_logic;
signal un2_cntr_c4 : std_logic;
signal \cntrZ0Z_0\ : std_logic;
signal \PWM_NUMZ0Z_0\ : std_logic;
signal un1_cntr_0 : std_logic;
signal \cntrZ0Z_5\ : std_logic;
signal \PWM_NUMZ0Z_5\ : std_logic;
signal \cntrZ0Z_6\ : std_logic;
signal \PORT1_c\ : std_logic;
signal \PORT_r3_1\ : std_logic;
signal \clk_div_RNI06L91Z0Z_11\ : std_logic;
signal clk_div_i_11 : std_logic;
signal \clk_divZ0Z_1\ : std_logic;
signal \clk_divZ0Z_0\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \clk_divZ0Z_2\ : std_logic;
signal clk_div_1_cry_1 : std_logic;
signal \clk_divZ0Z_3\ : std_logic;
signal clk_div_1_cry_2 : std_logic;
signal \clk_divZ0Z_4\ : std_logic;
signal clk_div_1_cry_3 : std_logic;
signal \clk_divZ0Z_5\ : std_logic;
signal clk_div_1_cry_4 : std_logic;
signal \clk_divZ0Z_6\ : std_logic;
signal clk_div_1_cry_5 : std_logic;
signal \clk_divZ0Z_7\ : std_logic;
signal clk_div_1_cry_6 : std_logic;
signal \clk_divZ0Z_8\ : std_logic;
signal clk_div_1_cry_7 : std_logic;
signal clk_div_1_cry_8 : std_logic;
signal \clk_divZ0Z_9\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal clk_div_1_cry_9 : std_logic;
signal \clk_divZ0Z_10\ : std_logic;
signal \CLK_0_c_g\ : std_logic;
signal \upZ0Z_2\ : std_logic;
signal \upZ0Z_1\ : std_logic;
signal \shift_ret_1_RNI69IQZ0\ : std_logic;
signal \BUT1_c\ : std_logic;
signal level_0 : std_logic;
signal \shift_0Z0Z_1\ : std_logic;
signal \upZ0Z_0\ : std_logic;
signal \shift_0Z0Z_2\ : std_logic;
signal \downZ0Z_1\ : std_logic;
signal \downZ0Z_2\ : std_logic;
signal \shift2_ret_1_RNITCIZ0Z51\ : std_logic;
signal level2_0 : std_logic;
signal \shift2_0Z0Z_1\ : std_logic;
signal \BUT2_c\ : std_logic;
signal \downZ0Z_0\ : std_logic;
signal un1_ten_ms_i : std_logic;
signal \shift2_0Z0Z_2\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \PORT1_wire\ : std_logic;
signal \BUT2_wire\ : std_logic;
signal \BUT1_wire\ : std_logic;

begin
    \CLK_wire\ <= CLK;
    PORT1 <= \PORT1_wire\;
    \BUT2_wire\ <= BUT2;
    \BUT1_wire\ <= BUT1;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__2678\,
            GLOBALBUFFEROUTPUT => \CLK_0_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2680\,
            DIN => \N__2679\,
            DOUT => \N__2678\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2680\,
            PADOUT => \N__2679\,
            PADIN => \N__2678\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORT1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2669\,
            DIN => \N__2668\,
            DOUT => \N__2667\,
            PACKAGEPIN => \PORT1_wire\
        );

    \PORT1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2669\,
            PADOUT => \N__2668\,
            PADIN => \N__2667\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1540\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUT2_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2660\,
            DIN => \N__2659\,
            DOUT => \N__2658\,
            PACKAGEPIN => \BUT2_wire\
        );

    \BUT2_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2660\,
            PADOUT => \N__2659\,
            PADIN => \N__2658\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BUT2_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUT1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2651\,
            DIN => \N__2650\,
            DOUT => \N__2649\,
            PACKAGEPIN => \BUT1_wire\
        );

    \BUT1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2651\,
            PADOUT => \N__2650\,
            PADIN => \N__2649\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BUT1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__597\ : CascadeMux
    port map (
            O => \N__2632\,
            I => \N__2628\
        );

    \I__596\ : InMux
    port map (
            O => \N__2631\,
            I => \N__2619\
        );

    \I__595\ : InMux
    port map (
            O => \N__2628\,
            I => \N__2619\
        );

    \I__594\ : InMux
    port map (
            O => \N__2627\,
            I => \N__2619\
        );

    \I__593\ : InMux
    port map (
            O => \N__2626\,
            I => \N__2616\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__2619\,
            I => \N__2613\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__2616\,
            I => \N__2610\
        );

    \I__590\ : Span4Mux_h
    port map (
            O => \N__2613\,
            I => \N__2607\
        );

    \I__589\ : Span4Mux_v
    port map (
            O => \N__2610\,
            I => \N__2604\
        );

    \I__588\ : Span4Mux_h
    port map (
            O => \N__2607\,
            I => \N__2601\
        );

    \I__587\ : Span4Mux_h
    port map (
            O => \N__2604\,
            I => \N__2598\
        );

    \I__586\ : Odrv4
    port map (
            O => \N__2601\,
            I => \BUT1_c\
        );

    \I__585\ : Odrv4
    port map (
            O => \N__2598\,
            I => \BUT1_c\
        );

    \I__584\ : CascadeMux
    port map (
            O => \N__2593\,
            I => \N__2589\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__2592\,
            I => \N__2586\
        );

    \I__582\ : InMux
    port map (
            O => \N__2589\,
            I => \N__2583\
        );

    \I__581\ : InMux
    port map (
            O => \N__2586\,
            I => \N__2580\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__2583\,
            I => level_0
        );

    \I__579\ : LocalMux
    port map (
            O => \N__2580\,
            I => level_0
        );

    \I__578\ : InMux
    port map (
            O => \N__2575\,
            I => \N__2570\
        );

    \I__577\ : InMux
    port map (
            O => \N__2574\,
            I => \N__2565\
        );

    \I__576\ : InMux
    port map (
            O => \N__2573\,
            I => \N__2565\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__2570\,
            I => \shift_0Z0Z_1\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__2565\,
            I => \shift_0Z0Z_1\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__2560\,
            I => \N__2555\
        );

    \I__572\ : InMux
    port map (
            O => \N__2559\,
            I => \N__2550\
        );

    \I__571\ : InMux
    port map (
            O => \N__2558\,
            I => \N__2550\
        );

    \I__570\ : InMux
    port map (
            O => \N__2555\,
            I => \N__2547\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__2550\,
            I => \N__2542\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__2547\,
            I => \N__2542\
        );

    \I__567\ : Span4Mux_v
    port map (
            O => \N__2542\,
            I => \N__2536\
        );

    \I__566\ : InMux
    port map (
            O => \N__2541\,
            I => \N__2531\
        );

    \I__565\ : InMux
    port map (
            O => \N__2540\,
            I => \N__2531\
        );

    \I__564\ : InMux
    port map (
            O => \N__2539\,
            I => \N__2528\
        );

    \I__563\ : Odrv4
    port map (
            O => \N__2536\,
            I => \upZ0Z_0\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__2531\,
            I => \upZ0Z_0\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__2528\,
            I => \upZ0Z_0\
        );

    \I__560\ : CEMux
    port map (
            O => \N__2521\,
            I => \N__2515\
        );

    \I__559\ : InMux
    port map (
            O => \N__2520\,
            I => \N__2508\
        );

    \I__558\ : InMux
    port map (
            O => \N__2519\,
            I => \N__2508\
        );

    \I__557\ : InMux
    port map (
            O => \N__2518\,
            I => \N__2508\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__2515\,
            I => \shift_0Z0Z_2\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__2508\,
            I => \shift_0Z0Z_2\
        );

    \I__554\ : InMux
    port map (
            O => \N__2503\,
            I => \N__2500\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__2500\,
            I => \N__2496\
        );

    \I__552\ : InMux
    port map (
            O => \N__2499\,
            I => \N__2493\
        );

    \I__551\ : Span4Mux_v
    port map (
            O => \N__2496\,
            I => \N__2488\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__2493\,
            I => \N__2485\
        );

    \I__549\ : InMux
    port map (
            O => \N__2492\,
            I => \N__2480\
        );

    \I__548\ : InMux
    port map (
            O => \N__2491\,
            I => \N__2480\
        );

    \I__547\ : Odrv4
    port map (
            O => \N__2488\,
            I => \downZ0Z_1\
        );

    \I__546\ : Odrv12
    port map (
            O => \N__2485\,
            I => \downZ0Z_1\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__2480\,
            I => \downZ0Z_1\
        );

    \I__544\ : InMux
    port map (
            O => \N__2473\,
            I => \N__2470\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__2470\,
            I => \N__2467\
        );

    \I__542\ : Span4Mux_v
    port map (
            O => \N__2467\,
            I => \N__2463\
        );

    \I__541\ : InMux
    port map (
            O => \N__2466\,
            I => \N__2460\
        );

    \I__540\ : Odrv4
    port map (
            O => \N__2463\,
            I => \downZ0Z_2\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__2460\,
            I => \downZ0Z_2\
        );

    \I__538\ : CEMux
    port map (
            O => \N__2455\,
            I => \N__2452\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__2452\,
            I => \N__2449\
        );

    \I__536\ : Span4Mux_v
    port map (
            O => \N__2449\,
            I => \N__2446\
        );

    \I__535\ : Span4Mux_s0_v
    port map (
            O => \N__2446\,
            I => \N__2443\
        );

    \I__534\ : Odrv4
    port map (
            O => \N__2443\,
            I => \shift2_ret_1_RNITCIZ0Z51\
        );

    \I__533\ : InMux
    port map (
            O => \N__2440\,
            I => \N__2436\
        );

    \I__532\ : InMux
    port map (
            O => \N__2439\,
            I => \N__2433\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__2436\,
            I => level2_0
        );

    \I__530\ : LocalMux
    port map (
            O => \N__2433\,
            I => level2_0
        );

    \I__529\ : CascadeMux
    port map (
            O => \N__2428\,
            I => \N__2424\
        );

    \I__528\ : InMux
    port map (
            O => \N__2427\,
            I => \N__2420\
        );

    \I__527\ : InMux
    port map (
            O => \N__2424\,
            I => \N__2415\
        );

    \I__526\ : InMux
    port map (
            O => \N__2423\,
            I => \N__2415\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__2420\,
            I => \shift2_0Z0Z_1\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__2415\,
            I => \shift2_0Z0Z_1\
        );

    \I__523\ : InMux
    port map (
            O => \N__2410\,
            I => \N__2406\
        );

    \I__522\ : CascadeMux
    port map (
            O => \N__2409\,
            I => \N__2402\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__2406\,
            I => \N__2398\
        );

    \I__520\ : InMux
    port map (
            O => \N__2405\,
            I => \N__2391\
        );

    \I__519\ : InMux
    port map (
            O => \N__2402\,
            I => \N__2391\
        );

    \I__518\ : InMux
    port map (
            O => \N__2401\,
            I => \N__2391\
        );

    \I__517\ : Span4Mux_v
    port map (
            O => \N__2398\,
            I => \N__2386\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__2391\,
            I => \N__2386\
        );

    \I__515\ : Span4Mux_h
    port map (
            O => \N__2386\,
            I => \N__2383\
        );

    \I__514\ : Odrv4
    port map (
            O => \N__2383\,
            I => \BUT2_c\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__2380\,
            I => \N__2377\
        );

    \I__512\ : InMux
    port map (
            O => \N__2377\,
            I => \N__2371\
        );

    \I__511\ : InMux
    port map (
            O => \N__2376\,
            I => \N__2371\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__2371\,
            I => \N__2366\
        );

    \I__509\ : InMux
    port map (
            O => \N__2370\,
            I => \N__2363\
        );

    \I__508\ : CascadeMux
    port map (
            O => \N__2369\,
            I => \N__2358\
        );

    \I__507\ : Span4Mux_v
    port map (
            O => \N__2366\,
            I => \N__2355\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__2363\,
            I => \N__2352\
        );

    \I__505\ : InMux
    port map (
            O => \N__2362\,
            I => \N__2347\
        );

    \I__504\ : InMux
    port map (
            O => \N__2361\,
            I => \N__2347\
        );

    \I__503\ : InMux
    port map (
            O => \N__2358\,
            I => \N__2344\
        );

    \I__502\ : Odrv4
    port map (
            O => \N__2355\,
            I => \downZ0Z_0\
        );

    \I__501\ : Odrv12
    port map (
            O => \N__2352\,
            I => \downZ0Z_0\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__2347\,
            I => \downZ0Z_0\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__2344\,
            I => \downZ0Z_0\
        );

    \I__498\ : ClkMux
    port map (
            O => \N__2335\,
            I => \N__2331\
        );

    \I__497\ : ClkMux
    port map (
            O => \N__2334\,
            I => \N__2327\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__2331\,
            I => \N__2322\
        );

    \I__495\ : ClkMux
    port map (
            O => \N__2330\,
            I => \N__2319\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__2327\,
            I => \N__2316\
        );

    \I__493\ : ClkMux
    port map (
            O => \N__2326\,
            I => \N__2313\
        );

    \I__492\ : ClkMux
    port map (
            O => \N__2325\,
            I => \N__2310\
        );

    \I__491\ : Span4Mux_s3_v
    port map (
            O => \N__2322\,
            I => \N__2306\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__2319\,
            I => \N__2303\
        );

    \I__489\ : Span4Mux_v
    port map (
            O => \N__2316\,
            I => \N__2298\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__2313\,
            I => \N__2298\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__2310\,
            I => \N__2295\
        );

    \I__486\ : ClkMux
    port map (
            O => \N__2309\,
            I => \N__2292\
        );

    \I__485\ : Span4Mux_h
    port map (
            O => \N__2306\,
            I => \N__2289\
        );

    \I__484\ : Span4Mux_v
    port map (
            O => \N__2303\,
            I => \N__2286\
        );

    \I__483\ : Span4Mux_h
    port map (
            O => \N__2298\,
            I => \N__2281\
        );

    \I__482\ : Span4Mux_h
    port map (
            O => \N__2295\,
            I => \N__2281\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__2292\,
            I => \N__2278\
        );

    \I__480\ : Odrv4
    port map (
            O => \N__2289\,
            I => un1_ten_ms_i
        );

    \I__479\ : Odrv4
    port map (
            O => \N__2286\,
            I => un1_ten_ms_i
        );

    \I__478\ : Odrv4
    port map (
            O => \N__2281\,
            I => un1_ten_ms_i
        );

    \I__477\ : Odrv12
    port map (
            O => \N__2278\,
            I => un1_ten_ms_i
        );

    \I__476\ : CEMux
    port map (
            O => \N__2269\,
            I => \N__2266\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__2266\,
            I => \N__2263\
        );

    \I__474\ : Sp12to4
    port map (
            O => \N__2263\,
            I => \N__2257\
        );

    \I__473\ : InMux
    port map (
            O => \N__2262\,
            I => \N__2250\
        );

    \I__472\ : InMux
    port map (
            O => \N__2261\,
            I => \N__2250\
        );

    \I__471\ : InMux
    port map (
            O => \N__2260\,
            I => \N__2250\
        );

    \I__470\ : Odrv12
    port map (
            O => \N__2257\,
            I => \shift2_0Z0Z_2\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__2250\,
            I => \shift2_0Z0Z_2\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__2245\,
            I => \N__2241\
        );

    \I__467\ : InMux
    port map (
            O => \N__2244\,
            I => \N__2238\
        );

    \I__466\ : InMux
    port map (
            O => \N__2241\,
            I => \N__2235\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__2238\,
            I => \clk_divZ0Z_8\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2235\,
            I => \clk_divZ0Z_8\
        );

    \I__463\ : InMux
    port map (
            O => \N__2230\,
            I => clk_div_1_cry_7
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__2227\,
            I => \N__2223\
        );

    \I__461\ : InMux
    port map (
            O => \N__2226\,
            I => \N__2220\
        );

    \I__460\ : InMux
    port map (
            O => \N__2223\,
            I => \N__2217\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__2220\,
            I => \clk_divZ0Z_9\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__2217\,
            I => \clk_divZ0Z_9\
        );

    \I__457\ : InMux
    port map (
            O => \N__2212\,
            I => \bfn_2_9_0_\
        );

    \I__456\ : InMux
    port map (
            O => \N__2209\,
            I => clk_div_1_cry_9
        );

    \I__455\ : InMux
    port map (
            O => \N__2206\,
            I => \N__2202\
        );

    \I__454\ : InMux
    port map (
            O => \N__2205\,
            I => \N__2199\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__2202\,
            I => \clk_divZ0Z_10\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__2199\,
            I => \clk_divZ0Z_10\
        );

    \I__451\ : ClkMux
    port map (
            O => \N__2194\,
            I => \N__2161\
        );

    \I__450\ : ClkMux
    port map (
            O => \N__2193\,
            I => \N__2161\
        );

    \I__449\ : ClkMux
    port map (
            O => \N__2192\,
            I => \N__2161\
        );

    \I__448\ : ClkMux
    port map (
            O => \N__2191\,
            I => \N__2161\
        );

    \I__447\ : ClkMux
    port map (
            O => \N__2190\,
            I => \N__2161\
        );

    \I__446\ : ClkMux
    port map (
            O => \N__2189\,
            I => \N__2161\
        );

    \I__445\ : ClkMux
    port map (
            O => \N__2188\,
            I => \N__2161\
        );

    \I__444\ : ClkMux
    port map (
            O => \N__2187\,
            I => \N__2161\
        );

    \I__443\ : ClkMux
    port map (
            O => \N__2186\,
            I => \N__2161\
        );

    \I__442\ : ClkMux
    port map (
            O => \N__2185\,
            I => \N__2161\
        );

    \I__441\ : ClkMux
    port map (
            O => \N__2184\,
            I => \N__2161\
        );

    \I__440\ : GlobalMux
    port map (
            O => \N__2161\,
            I => \N__2158\
        );

    \I__439\ : gio2CtrlBuf
    port map (
            O => \N__2158\,
            I => \CLK_0_c_g\
        );

    \I__438\ : InMux
    port map (
            O => \N__2155\,
            I => \N__2152\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__2152\,
            I => \N__2149\
        );

    \I__436\ : Span4Mux_s3_h
    port map (
            O => \N__2149\,
            I => \N__2145\
        );

    \I__435\ : InMux
    port map (
            O => \N__2148\,
            I => \N__2142\
        );

    \I__434\ : Odrv4
    port map (
            O => \N__2145\,
            I => \upZ0Z_2\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__2142\,
            I => \upZ0Z_2\
        );

    \I__432\ : InMux
    port map (
            O => \N__2137\,
            I => \N__2134\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2134\,
            I => \N__2130\
        );

    \I__430\ : InMux
    port map (
            O => \N__2133\,
            I => \N__2127\
        );

    \I__429\ : Span4Mux_v
    port map (
            O => \N__2130\,
            I => \N__2120\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2127\,
            I => \N__2120\
        );

    \I__427\ : InMux
    port map (
            O => \N__2126\,
            I => \N__2115\
        );

    \I__426\ : InMux
    port map (
            O => \N__2125\,
            I => \N__2115\
        );

    \I__425\ : Odrv4
    port map (
            O => \N__2120\,
            I => \upZ0Z_1\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__2115\,
            I => \upZ0Z_1\
        );

    \I__423\ : CEMux
    port map (
            O => \N__2110\,
            I => \N__2107\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2107\,
            I => \N__2104\
        );

    \I__421\ : Span4Mux_v
    port map (
            O => \N__2104\,
            I => \N__2101\
        );

    \I__420\ : Odrv4
    port map (
            O => \N__2101\,
            I => \shift_ret_1_RNI69IQZ0\
        );

    \I__419\ : InMux
    port map (
            O => \N__2098\,
            I => \N__2092\
        );

    \I__418\ : InMux
    port map (
            O => \N__2097\,
            I => \N__2087\
        );

    \I__417\ : InMux
    port map (
            O => \N__2096\,
            I => \N__2087\
        );

    \I__416\ : InMux
    port map (
            O => \N__2095\,
            I => \N__2084\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2092\,
            I => \N__2079\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__2087\,
            I => \N__2079\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__2084\,
            I => \clk_div_RNI06L91Z0Z_11\
        );

    \I__412\ : Odrv4
    port map (
            O => \N__2079\,
            I => \clk_div_RNI06L91Z0Z_11\
        );

    \I__411\ : InMux
    port map (
            O => \N__2074\,
            I => \N__2068\
        );

    \I__410\ : InMux
    port map (
            O => \N__2073\,
            I => \N__2063\
        );

    \I__409\ : InMux
    port map (
            O => \N__2072\,
            I => \N__2063\
        );

    \I__408\ : InMux
    port map (
            O => \N__2071\,
            I => \N__2060\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2068\,
            I => clk_div_i_11
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2063\,
            I => clk_div_i_11
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2060\,
            I => clk_div_i_11
        );

    \I__404\ : InMux
    port map (
            O => \N__2053\,
            I => \N__2048\
        );

    \I__403\ : InMux
    port map (
            O => \N__2052\,
            I => \N__2045\
        );

    \I__402\ : InMux
    port map (
            O => \N__2051\,
            I => \N__2042\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__2048\,
            I => \clk_divZ0Z_1\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__2045\,
            I => \clk_divZ0Z_1\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__2042\,
            I => \clk_divZ0Z_1\
        );

    \I__398\ : CascadeMux
    port map (
            O => \N__2035\,
            I => \N__2029\
        );

    \I__397\ : CascadeMux
    port map (
            O => \N__2034\,
            I => \N__2026\
        );

    \I__396\ : InMux
    port map (
            O => \N__2033\,
            I => \N__2023\
        );

    \I__395\ : InMux
    port map (
            O => \N__2032\,
            I => \N__2020\
        );

    \I__394\ : InMux
    port map (
            O => \N__2029\,
            I => \N__2017\
        );

    \I__393\ : InMux
    port map (
            O => \N__2026\,
            I => \N__2014\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__2023\,
            I => \clk_divZ0Z_0\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2020\,
            I => \clk_divZ0Z_0\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__2017\,
            I => \clk_divZ0Z_0\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__2014\,
            I => \clk_divZ0Z_0\
        );

    \I__388\ : CascadeMux
    port map (
            O => \N__2005\,
            I => \N__2001\
        );

    \I__387\ : InMux
    port map (
            O => \N__2004\,
            I => \N__1998\
        );

    \I__386\ : InMux
    port map (
            O => \N__2001\,
            I => \N__1995\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__1998\,
            I => \clk_divZ0Z_2\
        );

    \I__384\ : LocalMux
    port map (
            O => \N__1995\,
            I => \clk_divZ0Z_2\
        );

    \I__383\ : InMux
    port map (
            O => \N__1990\,
            I => clk_div_1_cry_1
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__1987\,
            I => \N__1983\
        );

    \I__381\ : InMux
    port map (
            O => \N__1986\,
            I => \N__1980\
        );

    \I__380\ : InMux
    port map (
            O => \N__1983\,
            I => \N__1977\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__1980\,
            I => \clk_divZ0Z_3\
        );

    \I__378\ : LocalMux
    port map (
            O => \N__1977\,
            I => \clk_divZ0Z_3\
        );

    \I__377\ : InMux
    port map (
            O => \N__1972\,
            I => clk_div_1_cry_2
        );

    \I__376\ : CascadeMux
    port map (
            O => \N__1969\,
            I => \N__1965\
        );

    \I__375\ : InMux
    port map (
            O => \N__1968\,
            I => \N__1962\
        );

    \I__374\ : InMux
    port map (
            O => \N__1965\,
            I => \N__1959\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__1962\,
            I => \clk_divZ0Z_4\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__1959\,
            I => \clk_divZ0Z_4\
        );

    \I__371\ : InMux
    port map (
            O => \N__1954\,
            I => clk_div_1_cry_3
        );

    \I__370\ : CascadeMux
    port map (
            O => \N__1951\,
            I => \N__1947\
        );

    \I__369\ : InMux
    port map (
            O => \N__1950\,
            I => \N__1944\
        );

    \I__368\ : InMux
    port map (
            O => \N__1947\,
            I => \N__1941\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__1944\,
            I => \clk_divZ0Z_5\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__1941\,
            I => \clk_divZ0Z_5\
        );

    \I__365\ : InMux
    port map (
            O => \N__1936\,
            I => clk_div_1_cry_4
        );

    \I__364\ : CascadeMux
    port map (
            O => \N__1933\,
            I => \N__1929\
        );

    \I__363\ : InMux
    port map (
            O => \N__1932\,
            I => \N__1926\
        );

    \I__362\ : InMux
    port map (
            O => \N__1929\,
            I => \N__1923\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__1926\,
            I => \clk_divZ0Z_6\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__1923\,
            I => \clk_divZ0Z_6\
        );

    \I__359\ : InMux
    port map (
            O => \N__1918\,
            I => clk_div_1_cry_5
        );

    \I__358\ : CascadeMux
    port map (
            O => \N__1915\,
            I => \N__1911\
        );

    \I__357\ : InMux
    port map (
            O => \N__1914\,
            I => \N__1908\
        );

    \I__356\ : InMux
    port map (
            O => \N__1911\,
            I => \N__1905\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__1908\,
            I => \clk_divZ0Z_7\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__1905\,
            I => \clk_divZ0Z_7\
        );

    \I__353\ : InMux
    port map (
            O => \N__1900\,
            I => clk_div_1_cry_6
        );

    \I__352\ : SRMux
    port map (
            O => \N__1897\,
            I => \N__1894\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__1894\,
            I => \N__1890\
        );

    \I__350\ : SRMux
    port map (
            O => \N__1893\,
            I => \N__1887\
        );

    \I__349\ : Span4Mux_s1_h
    port map (
            O => \N__1890\,
            I => \N__1882\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__1887\,
            I => \N__1882\
        );

    \I__347\ : Odrv4
    port map (
            O => \N__1882\,
            I => \PWM_NUM_RNIKTNT2Z0Z_0\
        );

    \I__346\ : CascadeMux
    port map (
            O => \N__1879\,
            I => \PWM_NUM_RNIKTNT2Z0Z_0_cascade_\
        );

    \I__345\ : CEMux
    port map (
            O => \N__1876\,
            I => \N__1873\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__1873\,
            I => \N_78_0\
        );

    \I__343\ : InMux
    port map (
            O => \N__1870\,
            I => \N__1866\
        );

    \I__342\ : InMux
    port map (
            O => \N__1869\,
            I => \N__1863\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__1866\,
            I => \PWM_NUMZ0Z_4\
        );

    \I__340\ : LocalMux
    port map (
            O => \N__1863\,
            I => \PWM_NUMZ0Z_4\
        );

    \I__339\ : InMux
    port map (
            O => \N__1858\,
            I => \N__1855\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__1855\,
            I => g0_3
        );

    \I__337\ : CascadeMux
    port map (
            O => \N__1852\,
            I => \N__1846\
        );

    \I__336\ : CascadeMux
    port map (
            O => \N__1851\,
            I => \N__1843\
        );

    \I__335\ : CascadeMux
    port map (
            O => \N__1850\,
            I => \N__1840\
        );

    \I__334\ : CascadeMux
    port map (
            O => \N__1849\,
            I => \N__1837\
        );

    \I__333\ : InMux
    port map (
            O => \N__1846\,
            I => \N__1833\
        );

    \I__332\ : InMux
    port map (
            O => \N__1843\,
            I => \N__1828\
        );

    \I__331\ : InMux
    port map (
            O => \N__1840\,
            I => \N__1828\
        );

    \I__330\ : InMux
    port map (
            O => \N__1837\,
            I => \N__1825\
        );

    \I__329\ : InMux
    port map (
            O => \N__1836\,
            I => \N__1822\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__1833\,
            I => \cntrZ0Z_4\
        );

    \I__327\ : LocalMux
    port map (
            O => \N__1828\,
            I => \cntrZ0Z_4\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__1825\,
            I => \cntrZ0Z_4\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__1822\,
            I => \cntrZ0Z_4\
        );

    \I__324\ : CEMux
    port map (
            O => \N__1813\,
            I => \N__1810\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__1810\,
            I => \N__1805\
        );

    \I__322\ : CEMux
    port map (
            O => \N__1809\,
            I => \N__1802\
        );

    \I__321\ : CEMux
    port map (
            O => \N__1808\,
            I => \N__1799\
        );

    \I__320\ : Span4Mux_v
    port map (
            O => \N__1805\,
            I => \N__1794\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__1802\,
            I => \N__1794\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__1799\,
            I => \N__1786\
        );

    \I__317\ : Span4Mux_h
    port map (
            O => \N__1794\,
            I => \N__1783\
        );

    \I__316\ : InMux
    port map (
            O => \N__1793\,
            I => \N__1774\
        );

    \I__315\ : InMux
    port map (
            O => \N__1792\,
            I => \N__1774\
        );

    \I__314\ : InMux
    port map (
            O => \N__1791\,
            I => \N__1774\
        );

    \I__313\ : InMux
    port map (
            O => \N__1790\,
            I => \N__1774\
        );

    \I__312\ : InMux
    port map (
            O => \N__1789\,
            I => \N__1771\
        );

    \I__311\ : Odrv4
    port map (
            O => \N__1786\,
            I => \clk_div_RNIM1KP1Z0Z_11\
        );

    \I__310\ : Odrv4
    port map (
            O => \N__1783\,
            I => \clk_div_RNIM1KP1Z0Z_11\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__1774\,
            I => \clk_div_RNIM1KP1Z0Z_11\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__1771\,
            I => \clk_div_RNIM1KP1Z0Z_11\
        );

    \I__307\ : InMux
    port map (
            O => \N__1762\,
            I => \N__1758\
        );

    \I__306\ : InMux
    port map (
            O => \N__1761\,
            I => \N__1753\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__1758\,
            I => \N__1750\
        );

    \I__304\ : InMux
    port map (
            O => \N__1757\,
            I => \N__1745\
        );

    \I__303\ : InMux
    port map (
            O => \N__1756\,
            I => \N__1745\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__1753\,
            I => \cntrZ0Z_3\
        );

    \I__301\ : Odrv4
    port map (
            O => \N__1750\,
            I => \cntrZ0Z_3\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__1745\,
            I => \cntrZ0Z_3\
        );

    \I__299\ : InMux
    port map (
            O => \N__1738\,
            I => \N__1732\
        );

    \I__298\ : InMux
    port map (
            O => \N__1737\,
            I => \N__1729\
        );

    \I__297\ : InMux
    port map (
            O => \N__1736\,
            I => \N__1726\
        );

    \I__296\ : InMux
    port map (
            O => \N__1735\,
            I => \N__1723\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__1732\,
            I => \cntrZ0Z_2\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__1729\,
            I => \cntrZ0Z_2\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__1726\,
            I => \cntrZ0Z_2\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__1723\,
            I => \cntrZ0Z_2\
        );

    \I__291\ : InMux
    port map (
            O => \N__1714\,
            I => \N__1707\
        );

    \I__290\ : InMux
    port map (
            O => \N__1713\,
            I => \N__1702\
        );

    \I__289\ : InMux
    port map (
            O => \N__1712\,
            I => \N__1702\
        );

    \I__288\ : InMux
    port map (
            O => \N__1711\,
            I => \N__1699\
        );

    \I__287\ : InMux
    port map (
            O => \N__1710\,
            I => \N__1696\
        );

    \I__286\ : LocalMux
    port map (
            O => \N__1707\,
            I => \cntrZ0Z_1\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__1702\,
            I => \cntrZ0Z_1\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__1699\,
            I => \cntrZ0Z_1\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__1696\,
            I => \cntrZ0Z_1\
        );

    \I__282\ : InMux
    port map (
            O => \N__1687\,
            I => \N__1682\
        );

    \I__281\ : InMux
    port map (
            O => \N__1686\,
            I => \N__1677\
        );

    \I__280\ : InMux
    port map (
            O => \N__1685\,
            I => \N__1677\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__1682\,
            I => un2_cntr_c4
        );

    \I__278\ : LocalMux
    port map (
            O => \N__1677\,
            I => un2_cntr_c4
        );

    \I__277\ : CascadeMux
    port map (
            O => \N__1672\,
            I => \N__1665\
        );

    \I__276\ : CascadeMux
    port map (
            O => \N__1671\,
            I => \N__1662\
        );

    \I__275\ : CascadeMux
    port map (
            O => \N__1670\,
            I => \N__1657\
        );

    \I__274\ : CascadeMux
    port map (
            O => \N__1669\,
            I => \N__1654\
        );

    \I__273\ : InMux
    port map (
            O => \N__1668\,
            I => \N__1651\
        );

    \I__272\ : InMux
    port map (
            O => \N__1665\,
            I => \N__1648\
        );

    \I__271\ : InMux
    port map (
            O => \N__1662\,
            I => \N__1643\
        );

    \I__270\ : InMux
    port map (
            O => \N__1661\,
            I => \N__1643\
        );

    \I__269\ : InMux
    port map (
            O => \N__1660\,
            I => \N__1638\
        );

    \I__268\ : InMux
    port map (
            O => \N__1657\,
            I => \N__1638\
        );

    \I__267\ : InMux
    port map (
            O => \N__1654\,
            I => \N__1635\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__1651\,
            I => \cntrZ0Z_0\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__1648\,
            I => \cntrZ0Z_0\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__1643\,
            I => \cntrZ0Z_0\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__1638\,
            I => \cntrZ0Z_0\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__1635\,
            I => \cntrZ0Z_0\
        );

    \I__261\ : InMux
    port map (
            O => \N__1624\,
            I => \N__1620\
        );

    \I__260\ : InMux
    port map (
            O => \N__1623\,
            I => \N__1617\
        );

    \I__259\ : LocalMux
    port map (
            O => \N__1620\,
            I => \N__1612\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__1617\,
            I => \N__1612\
        );

    \I__257\ : Odrv4
    port map (
            O => \N__1612\,
            I => \PWM_NUMZ0Z_0\
        );

    \I__256\ : InMux
    port map (
            O => \N__1609\,
            I => \N__1606\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__1606\,
            I => un1_cntr_0
        );

    \I__254\ : CascadeMux
    port map (
            O => \N__1603\,
            I => \N__1597\
        );

    \I__253\ : InMux
    port map (
            O => \N__1602\,
            I => \N__1594\
        );

    \I__252\ : InMux
    port map (
            O => \N__1601\,
            I => \N__1591\
        );

    \I__251\ : InMux
    port map (
            O => \N__1600\,
            I => \N__1588\
        );

    \I__250\ : InMux
    port map (
            O => \N__1597\,
            I => \N__1585\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__1594\,
            I => \cntrZ0Z_5\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__1591\,
            I => \cntrZ0Z_5\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__1588\,
            I => \cntrZ0Z_5\
        );

    \I__246\ : LocalMux
    port map (
            O => \N__1585\,
            I => \cntrZ0Z_5\
        );

    \I__245\ : InMux
    port map (
            O => \N__1576\,
            I => \N__1573\
        );

    \I__244\ : LocalMux
    port map (
            O => \N__1573\,
            I => \N__1569\
        );

    \I__243\ : InMux
    port map (
            O => \N__1572\,
            I => \N__1566\
        );

    \I__242\ : Odrv4
    port map (
            O => \N__1569\,
            I => \PWM_NUMZ0Z_5\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__1566\,
            I => \PWM_NUMZ0Z_5\
        );

    \I__240\ : CascadeMux
    port map (
            O => \N__1561\,
            I => \N__1557\
        );

    \I__239\ : CascadeMux
    port map (
            O => \N__1560\,
            I => \N__1553\
        );

    \I__238\ : InMux
    port map (
            O => \N__1557\,
            I => \N__1550\
        );

    \I__237\ : InMux
    port map (
            O => \N__1556\,
            I => \N__1545\
        );

    \I__236\ : InMux
    port map (
            O => \N__1553\,
            I => \N__1545\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__1550\,
            I => \cntrZ0Z_6\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__1545\,
            I => \cntrZ0Z_6\
        );

    \I__233\ : IoInMux
    port map (
            O => \N__1540\,
            I => \N__1537\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__1537\,
            I => \N__1534\
        );

    \I__231\ : Span12Mux_s1_h
    port map (
            O => \N__1534\,
            I => \N__1529\
        );

    \I__230\ : InMux
    port map (
            O => \N__1533\,
            I => \N__1526\
        );

    \I__229\ : InMux
    port map (
            O => \N__1532\,
            I => \N__1523\
        );

    \I__228\ : Odrv12
    port map (
            O => \N__1529\,
            I => \PORT1_c\
        );

    \I__227\ : LocalMux
    port map (
            O => \N__1526\,
            I => \PORT1_c\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__1523\,
            I => \PORT1_c\
        );

    \I__225\ : CascadeMux
    port map (
            O => \N__1516\,
            I => \N__1513\
        );

    \I__224\ : InMux
    port map (
            O => \N__1513\,
            I => \N__1510\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__1510\,
            I => \N__1507\
        );

    \I__222\ : Odrv4
    port map (
            O => \N__1507\,
            I => \PORT_r3_1\
        );

    \I__221\ : InMux
    port map (
            O => \N__1504\,
            I => \N__1498\
        );

    \I__220\ : InMux
    port map (
            O => \N__1503\,
            I => \N__1498\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__1498\,
            I => \PWM_NUMZ0Z_3\
        );

    \I__218\ : CascadeMux
    port map (
            O => \N__1495\,
            I => \N__1492\
        );

    \I__217\ : InMux
    port map (
            O => \N__1492\,
            I => \N__1489\
        );

    \I__216\ : LocalMux
    port map (
            O => \N__1489\,
            I => \PWM_NUMZ0Z_1\
        );

    \I__215\ : InMux
    port map (
            O => \N__1486\,
            I => \N__1473\
        );

    \I__214\ : InMux
    port map (
            O => \N__1485\,
            I => \N__1473\
        );

    \I__213\ : InMux
    port map (
            O => \N__1484\,
            I => \N__1473\
        );

    \I__212\ : InMux
    port map (
            O => \N__1483\,
            I => \N__1473\
        );

    \I__211\ : InMux
    port map (
            O => \N__1482\,
            I => \N__1470\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__1473\,
            I => \howZ0Z_0\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__1470\,
            I => \howZ0Z_0\
        );

    \I__208\ : InMux
    port map (
            O => \N__1465\,
            I => \N__1449\
        );

    \I__207\ : InMux
    port map (
            O => \N__1464\,
            I => \N__1449\
        );

    \I__206\ : InMux
    port map (
            O => \N__1463\,
            I => \N__1449\
        );

    \I__205\ : InMux
    port map (
            O => \N__1462\,
            I => \N__1449\
        );

    \I__204\ : InMux
    port map (
            O => \N__1461\,
            I => \N__1449\
        );

    \I__203\ : InMux
    port map (
            O => \N__1460\,
            I => \N__1446\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__1449\,
            I => \howZ0Z_2\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__1446\,
            I => \howZ0Z_2\
        );

    \I__200\ : InMux
    port map (
            O => \N__1441\,
            I => \N__1428\
        );

    \I__199\ : InMux
    port map (
            O => \N__1440\,
            I => \N__1428\
        );

    \I__198\ : InMux
    port map (
            O => \N__1439\,
            I => \N__1428\
        );

    \I__197\ : InMux
    port map (
            O => \N__1438\,
            I => \N__1428\
        );

    \I__196\ : InMux
    port map (
            O => \N__1437\,
            I => \N__1425\
        );

    \I__195\ : LocalMux
    port map (
            O => \N__1428\,
            I => \howZ0Z_1\
        );

    \I__194\ : LocalMux
    port map (
            O => \N__1425\,
            I => \howZ0Z_1\
        );

    \I__193\ : InMux
    port map (
            O => \N__1420\,
            I => \N__1417\
        );

    \I__192\ : LocalMux
    port map (
            O => \N__1417\,
            I => \PWM_NUMZ0Z_2\
        );

    \I__191\ : InMux
    port map (
            O => \N__1414\,
            I => \N__1411\
        );

    \I__190\ : LocalMux
    port map (
            O => \N__1411\,
            I => \PORT_r3_2\
        );

    \I__189\ : InMux
    port map (
            O => \N__1408\,
            I => \N__1402\
        );

    \I__188\ : InMux
    port map (
            O => \N__1407\,
            I => \N__1402\
        );

    \I__187\ : LocalMux
    port map (
            O => \N__1402\,
            I => \PORT_r3_3\
        );

    \I__186\ : InMux
    port map (
            O => \N__1399\,
            I => \N__1396\
        );

    \I__185\ : LocalMux
    port map (
            O => \N__1396\,
            I => g0_2
        );

    \I__184\ : CascadeMux
    port map (
            O => \N__1393\,
            I => \g0_4_cascade_\
        );

    \I__183\ : InMux
    port map (
            O => \N__1390\,
            I => \N__1386\
        );

    \I__182\ : InMux
    port map (
            O => \N__1389\,
            I => \N__1383\
        );

    \I__181\ : LocalMux
    port map (
            O => \N__1386\,
            I => \delayZ0Z_10\
        );

    \I__180\ : LocalMux
    port map (
            O => \N__1383\,
            I => \delayZ0Z_10\
        );

    \I__179\ : CascadeMux
    port map (
            O => \N__1378\,
            I => \N__1375\
        );

    \I__178\ : InMux
    port map (
            O => \N__1375\,
            I => \N__1371\
        );

    \I__177\ : InMux
    port map (
            O => \N__1374\,
            I => \N__1368\
        );

    \I__176\ : LocalMux
    port map (
            O => \N__1371\,
            I => \delayZ0Z_8\
        );

    \I__175\ : LocalMux
    port map (
            O => \N__1368\,
            I => \delayZ0Z_8\
        );

    \I__174\ : InMux
    port map (
            O => \N__1363\,
            I => \N__1359\
        );

    \I__173\ : InMux
    port map (
            O => \N__1362\,
            I => \N__1356\
        );

    \I__172\ : LocalMux
    port map (
            O => \N__1359\,
            I => \delayZ0Z_9\
        );

    \I__171\ : LocalMux
    port map (
            O => \N__1356\,
            I => \delayZ0Z_9\
        );

    \I__170\ : InMux
    port map (
            O => \N__1351\,
            I => \N__1347\
        );

    \I__169\ : InMux
    port map (
            O => \N__1350\,
            I => \N__1344\
        );

    \I__168\ : LocalMux
    port map (
            O => \N__1347\,
            I => \delayZ0Z_0\
        );

    \I__167\ : LocalMux
    port map (
            O => \N__1344\,
            I => \delayZ0Z_0\
        );

    \I__166\ : InMux
    port map (
            O => \N__1339\,
            I => \N__1335\
        );

    \I__165\ : InMux
    port map (
            O => \N__1338\,
            I => \N__1332\
        );

    \I__164\ : LocalMux
    port map (
            O => \N__1335\,
            I => \delayZ0Z_3\
        );

    \I__163\ : LocalMux
    port map (
            O => \N__1332\,
            I => \delayZ0Z_3\
        );

    \I__162\ : CascadeMux
    port map (
            O => \N__1327\,
            I => \N__1324\
        );

    \I__161\ : InMux
    port map (
            O => \N__1324\,
            I => \N__1320\
        );

    \I__160\ : InMux
    port map (
            O => \N__1323\,
            I => \N__1317\
        );

    \I__159\ : LocalMux
    port map (
            O => \N__1320\,
            I => \delayZ0Z_1\
        );

    \I__158\ : LocalMux
    port map (
            O => \N__1317\,
            I => \delayZ0Z_1\
        );

    \I__157\ : InMux
    port map (
            O => \N__1312\,
            I => \N__1308\
        );

    \I__156\ : InMux
    port map (
            O => \N__1311\,
            I => \N__1305\
        );

    \I__155\ : LocalMux
    port map (
            O => \N__1308\,
            I => \delayZ0Z_2\
        );

    \I__154\ : LocalMux
    port map (
            O => \N__1305\,
            I => \delayZ0Z_2\
        );

    \I__153\ : InMux
    port map (
            O => \N__1300\,
            I => \N__1297\
        );

    \I__152\ : LocalMux
    port map (
            O => \N__1297\,
            I => un1_ten_ms_7
        );

    \I__151\ : InMux
    port map (
            O => \N__1294\,
            I => \N__1291\
        );

    \I__150\ : LocalMux
    port map (
            O => \N__1291\,
            I => un1_ten_ms_9
        );

    \I__149\ : CascadeMux
    port map (
            O => \N__1288\,
            I => \un1_ten_ms_8_cascade_\
        );

    \I__148\ : InMux
    port map (
            O => \N__1285\,
            I => \N__1282\
        );

    \I__147\ : LocalMux
    port map (
            O => \N__1282\,
            I => un1_ten_ms_10
        );

    \I__146\ : InMux
    port map (
            O => \N__1279\,
            I => \N__1276\
        );

    \I__145\ : LocalMux
    port map (
            O => \N__1276\,
            I => how_1_c2
        );

    \I__144\ : InMux
    port map (
            O => \N__1273\,
            I => clk_div_2_cry_10
        );

    \I__143\ : InMux
    port map (
            O => \N__1270\,
            I => \N__1266\
        );

    \I__142\ : InMux
    port map (
            O => \N__1269\,
            I => \N__1263\
        );

    \I__141\ : LocalMux
    port map (
            O => \N__1266\,
            I => \delayZ0Z_6\
        );

    \I__140\ : LocalMux
    port map (
            O => \N__1263\,
            I => \delayZ0Z_6\
        );

    \I__139\ : InMux
    port map (
            O => \N__1258\,
            I => \N__1254\
        );

    \I__138\ : InMux
    port map (
            O => \N__1257\,
            I => \N__1251\
        );

    \I__137\ : LocalMux
    port map (
            O => \N__1254\,
            I => \delayZ0Z_5\
        );

    \I__136\ : LocalMux
    port map (
            O => \N__1251\,
            I => \delayZ0Z_5\
        );

    \I__135\ : InMux
    port map (
            O => \N__1246\,
            I => \N__1242\
        );

    \I__134\ : InMux
    port map (
            O => \N__1245\,
            I => \N__1239\
        );

    \I__133\ : LocalMux
    port map (
            O => \N__1242\,
            I => \delayZ0Z_4\
        );

    \I__132\ : LocalMux
    port map (
            O => \N__1239\,
            I => \delayZ0Z_4\
        );

    \I__131\ : InMux
    port map (
            O => \N__1234\,
            I => \N__1230\
        );

    \I__130\ : InMux
    port map (
            O => \N__1233\,
            I => \N__1227\
        );

    \I__129\ : LocalMux
    port map (
            O => \N__1230\,
            I => \delayZ0Z_7\
        );

    \I__128\ : LocalMux
    port map (
            O => \N__1227\,
            I => \delayZ0Z_7\
        );

    \I__127\ : InMux
    port map (
            O => \N__1222\,
            I => \bfn_1_3_0_\
        );

    \I__126\ : InMux
    port map (
            O => \N__1219\,
            I => delay_cry_8
        );

    \I__125\ : InMux
    port map (
            O => \N__1216\,
            I => delay_cry_9
        );

    \I__124\ : InMux
    port map (
            O => \N__1213\,
            I => delay_cry_10
        );

    \I__123\ : InMux
    port map (
            O => \N__1210\,
            I => delay_cry_11
        );

    \I__122\ : InMux
    port map (
            O => \N__1207\,
            I => delay_cry_12
        );

    \I__121\ : InMux
    port map (
            O => \N__1204\,
            I => delay_cry_13
        );

    \I__120\ : InMux
    port map (
            O => \N__1201\,
            I => \N__1195\
        );

    \I__119\ : InMux
    port map (
            O => \N__1200\,
            I => \N__1195\
        );

    \I__118\ : LocalMux
    port map (
            O => \N__1195\,
            I => \delayZ0Z_14\
        );

    \I__117\ : InMux
    port map (
            O => \N__1192\,
            I => \N__1186\
        );

    \I__116\ : InMux
    port map (
            O => \N__1191\,
            I => \N__1186\
        );

    \I__115\ : LocalMux
    port map (
            O => \N__1186\,
            I => \delayZ0Z_13\
        );

    \I__114\ : CascadeMux
    port map (
            O => \N__1183\,
            I => \N__1180\
        );

    \I__113\ : InMux
    port map (
            O => \N__1180\,
            I => \N__1174\
        );

    \I__112\ : InMux
    port map (
            O => \N__1179\,
            I => \N__1174\
        );

    \I__111\ : LocalMux
    port map (
            O => \N__1174\,
            I => \delayZ0Z_12\
        );

    \I__110\ : InMux
    port map (
            O => \N__1171\,
            I => \N__1165\
        );

    \I__109\ : InMux
    port map (
            O => \N__1170\,
            I => \N__1165\
        );

    \I__108\ : LocalMux
    port map (
            O => \N__1165\,
            I => \delayZ0Z_11\
        );

    \I__107\ : InMux
    port map (
            O => \N__1162\,
            I => \bfn_1_2_0_\
        );

    \I__106\ : InMux
    port map (
            O => \N__1159\,
            I => delay_cry_0
        );

    \I__105\ : InMux
    port map (
            O => \N__1156\,
            I => delay_cry_1
        );

    \I__104\ : InMux
    port map (
            O => \N__1153\,
            I => delay_cry_2
        );

    \I__103\ : InMux
    port map (
            O => \N__1150\,
            I => delay_cry_3
        );

    \I__102\ : InMux
    port map (
            O => \N__1147\,
            I => delay_cry_4
        );

    \I__101\ : InMux
    port map (
            O => \N__1144\,
            I => delay_cry_5
        );

    \I__100\ : InMux
    port map (
            O => \N__1141\,
            I => delay_cry_6
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => clk_div_2_cry_8,
            carryinitout => \bfn_1_8_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => clk_div_1_cry_8,
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_1_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_2_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => delay_cry_7,
            carryinitout => \bfn_1_3_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \delay_0_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1350\,
            in2 => \_gnd_net_\,
            in3 => \N__1162\,
            lcout => \delayZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_2_0_\,
            carryout => delay_cry_0,
            clk => \N__2194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_1_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1323\,
            in2 => \_gnd_net_\,
            in3 => \N__1159\,
            lcout => \delayZ0Z_1\,
            ltout => OPEN,
            carryin => delay_cry_0,
            carryout => delay_cry_1,
            clk => \N__2194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_2_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1311\,
            in2 => \_gnd_net_\,
            in3 => \N__1156\,
            lcout => \delayZ0Z_2\,
            ltout => OPEN,
            carryin => delay_cry_1,
            carryout => delay_cry_2,
            clk => \N__2194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_3_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1338\,
            in2 => \_gnd_net_\,
            in3 => \N__1153\,
            lcout => \delayZ0Z_3\,
            ltout => OPEN,
            carryin => delay_cry_2,
            carryout => delay_cry_3,
            clk => \N__2194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_4_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1245\,
            in2 => \_gnd_net_\,
            in3 => \N__1150\,
            lcout => \delayZ0Z_4\,
            ltout => OPEN,
            carryin => delay_cry_3,
            carryout => delay_cry_4,
            clk => \N__2194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_5_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1257\,
            in2 => \_gnd_net_\,
            in3 => \N__1147\,
            lcout => \delayZ0Z_5\,
            ltout => OPEN,
            carryin => delay_cry_4,
            carryout => delay_cry_5,
            clk => \N__2194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_6_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1269\,
            in2 => \_gnd_net_\,
            in3 => \N__1144\,
            lcout => \delayZ0Z_6\,
            ltout => OPEN,
            carryin => delay_cry_5,
            carryout => delay_cry_6,
            clk => \N__2194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_7_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1233\,
            in2 => \_gnd_net_\,
            in3 => \N__1141\,
            lcout => \delayZ0Z_7\,
            ltout => OPEN,
            carryin => delay_cry_6,
            carryout => delay_cry_7,
            clk => \N__2194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_8_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1374\,
            in2 => \_gnd_net_\,
            in3 => \N__1222\,
            lcout => \delayZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => delay_cry_8,
            clk => \N__2192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_9_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1362\,
            in2 => \_gnd_net_\,
            in3 => \N__1219\,
            lcout => \delayZ0Z_9\,
            ltout => OPEN,
            carryin => delay_cry_8,
            carryout => delay_cry_9,
            clk => \N__2192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_10_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1389\,
            in2 => \_gnd_net_\,
            in3 => \N__1216\,
            lcout => \delayZ0Z_10\,
            ltout => OPEN,
            carryin => delay_cry_9,
            carryout => delay_cry_10,
            clk => \N__2192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_11_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1170\,
            in2 => \_gnd_net_\,
            in3 => \N__1213\,
            lcout => \delayZ0Z_11\,
            ltout => OPEN,
            carryin => delay_cry_10,
            carryout => delay_cry_11,
            clk => \N__2192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_12_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1179\,
            in2 => \_gnd_net_\,
            in3 => \N__1210\,
            lcout => \delayZ0Z_12\,
            ltout => OPEN,
            carryin => delay_cry_11,
            carryout => delay_cry_12,
            clk => \N__2192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_13_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1191\,
            in2 => \_gnd_net_\,
            in3 => \N__1207\,
            lcout => \delayZ0Z_13\,
            ltout => OPEN,
            carryin => delay_cry_12,
            carryout => delay_cry_13,
            clk => \N__2192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_14_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1200\,
            in2 => \_gnd_net_\,
            in3 => \N__1204\,
            lcout => \delayZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2192\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_RNIABQR_14_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1201\,
            in1 => \N__1192\,
            in2 => \N__1183\,
            in3 => \N__1171\,
            lcout => un1_ten_ms_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_esr_3_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__1761\,
            in1 => \N__1738\,
            in2 => \N__1672\,
            in3 => \N__1714\,
            lcout => \cntrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2189\,
            ce => \N__1876\,
            sr => \N__1897\
        );

    \cntr_2_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__1737\,
            in1 => \N__1713\,
            in2 => \N__1671\,
            in3 => \N__1792\,
            lcout => \cntrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2186\,
            ce => 'H',
            sr => \N__1893\
        );

    \cntr_4_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100001111000"
        )
    port map (
            in0 => \N__1791\,
            in1 => \N__1685\,
            in2 => \N__1851\,
            in3 => \_gnd_net_\,
            lcout => \cntrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2186\,
            ce => 'H',
            sr => \N__1893\
        );

    \cntr_5_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__1793\,
            in1 => \N__1601\,
            in2 => \N__1850\,
            in3 => \N__1686\,
            lcout => \cntrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2186\,
            ce => 'H',
            sr => \N__1893\
        );

    \cntr_1_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__1661\,
            in1 => \N__1712\,
            in2 => \_gnd_net_\,
            in3 => \N__1790\,
            lcout => \cntrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2186\,
            ce => 'H',
            sr => \N__1893\
        );

    \cntr_0_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__1668\,
            in1 => \N__2074\,
            in2 => \_gnd_net_\,
            in3 => \N__2098\,
            lcout => \cntrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2186\,
            ce => 'H',
            sr => \N__1893\
        );

    \clk_div_RNI91U1_1_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2051\,
            in2 => \N__2034\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => clk_div_2_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIF3T2_2_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2005\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_1,
            carryout => clk_div_2_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIM6S3_3_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1987\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_2,
            carryout => clk_div_2_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIUAR4_4_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1969\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_3,
            carryout => clk_div_2_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNI7GQ5_5_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1951\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_4,
            carryout => clk_div_2_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIHMP6_6_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1933\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_5,
            carryout => clk_div_2_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNISTO7_7_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1915\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_6,
            carryout => clk_div_2_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNI86O8_8_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2245\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_7,
            carryout => clk_div_2_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNILFN9_9_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2227\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_8_0_\,
            carryout => clk_div_2_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIAAMP_10_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2205\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_9,
            carryout => clk_div_2_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNI06L91_11_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2071\,
            in2 => \_gnd_net_\,
            in3 => \N__1273\,
            lcout => \clk_div_RNI06L91Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_1_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2033\,
            in2 => \_gnd_net_\,
            in3 => \N__2053\,
            lcout => \clk_divZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_RNIKNK01_4_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__1270\,
            in1 => \N__1258\,
            in2 => \_gnd_net_\,
            in3 => \N__1246\,
            lcout => un1_ten_ms_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_RNI5HJ71_10_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1234\,
            in1 => \N__1390\,
            in2 => \N__1378\,
            in3 => \N__1363\,
            lcout => un1_ten_ms_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_RNI2HGB1_0_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__1351\,
            in1 => \N__1339\,
            in2 => \N__1327\,
            in3 => \N__1312\,
            lcout => OPEN,
            ltout => \un1_ten_ms_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \delay_RNI55JF4_10_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1300\,
            in1 => \N__1294\,
            in2 => \N__1288\,
            in3 => \N__1285\,
            lcout => un1_ten_ms_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \how_RNO_0_2_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001010111011"
        )
    port map (
            in0 => \N__2133\,
            in1 => \N__2499\,
            in2 => \N__2560\,
            in3 => \N__2370\,
            lcout => how_1_c2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \how_1_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110001110011100"
        )
    port map (
            in0 => \N__2559\,
            in1 => \N__2137\,
            in2 => \N__2380\,
            in3 => \N__2503\,
            lcout => \howZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2193\,
            ce => \N__1808\,
            sr => \_gnd_net_\
        );

    \how_0_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2558\,
            in2 => \_gnd_net_\,
            in3 => \N__2376\,
            lcout => \howZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2193\,
            ce => \N__1808\,
            sr => \_gnd_net_\
        );

    \PWM_NUM_0_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1460\,
            in2 => \_gnd_net_\,
            in3 => \N__1482\,
            lcout => \PWM_NUMZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2193\,
            ce => \N__1808\,
            sr => \_gnd_net_\
        );

    \how_2_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010011001"
        )
    port map (
            in0 => \N__1279\,
            in1 => \N__2155\,
            in2 => \_gnd_net_\,
            in3 => \N__2473\,
            lcout => \howZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2193\,
            ce => \N__1808\,
            sr => \_gnd_net_\
        );

    \PORT_r_RNO_1_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__1757\,
            in1 => \N__1870\,
            in2 => \N__1849\,
            in3 => \N__1504\,
            lcout => \PORT_r3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM_NUM_3_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__1485\,
            in1 => \N__1464\,
            in2 => \_gnd_net_\,
            in3 => \N__1440\,
            lcout => \PWM_NUMZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2191\,
            ce => \N__1813\,
            sr => \_gnd_net_\
        );

    \PWM_NUM_RNIDRQK_3_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__1756\,
            in1 => \N__1572\,
            in2 => \N__1603\,
            in3 => \N__1503\,
            lcout => g0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM_NUM_5_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__1486\,
            in1 => \N__1465\,
            in2 => \_gnd_net_\,
            in3 => \N__1441\,
            lcout => \PWM_NUMZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2191\,
            ce => \N__1813\,
            sr => \_gnd_net_\
        );

    \PWM_NUM_4_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__1461\,
            in1 => \N__1437\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PWM_NUMZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2191\,
            ce => \N__1813\,
            sr => \_gnd_net_\
        );

    \PWM_NUM_1_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101100110"
        )
    port map (
            in0 => \N__1483\,
            in1 => \N__1462\,
            in2 => \_gnd_net_\,
            in3 => \N__1438\,
            lcout => \PWM_NUMZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2191\,
            ce => \N__1813\,
            sr => \_gnd_net_\
        );

    \PWM_NUM_RNIQIR6_1_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__1735\,
            in1 => \N__1710\,
            in2 => \N__1495\,
            in3 => \N__1420\,
            lcout => \PORT_r3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM_NUM_2_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001000100"
        )
    port map (
            in0 => \N__1484\,
            in1 => \N__1463\,
            in2 => \_gnd_net_\,
            in3 => \N__1439\,
            lcout => \PWM_NUMZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2191\,
            ce => \N__1813\,
            sr => \_gnd_net_\
        );

    \PORT_r_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__1408\,
            in1 => \N__1414\,
            in2 => \N__1516\,
            in3 => \N__1609\,
            lcout => \PORT1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2190\,
            ce => \N__1809\,
            sr => \_gnd_net_\
        );

    \PWM_NUM_RNIQ48Q_0_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000100000000"
        )
    port map (
            in0 => \N__1623\,
            in1 => \N__2072\,
            in2 => \N__1669\,
            in3 => \N__1407\,
            lcout => OPEN,
            ltout => \g0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM_NUM_RNIKTNT2_0_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1858\,
            in1 => \N__1399\,
            in2 => \N__1393\,
            in3 => \N__2097\,
            lcout => \PWM_NUM_RNIKTNT2Z0Z_0\,
            ltout => \PWM_NUM_RNIKTNT2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_esr_RNO_0_3_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1879\,
            in3 => \N__1789\,
            lcout => \N_78_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIM1KP1_11_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__2073\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2096\,
            lcout => \clk_div_RNIM1KP1Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PWM_NUM_RNIDNV4_4_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001001"
        )
    port map (
            in0 => \N__1869\,
            in1 => \N__1836\,
            in2 => \N__1560\,
            in3 => \N__1532\,
            lcout => g0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_6_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__1556\,
            in1 => \N__1687\,
            in2 => \N__1852\,
            in3 => \N__1602\,
            lcout => \cntrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2190\,
            ce => \N__1809\,
            sr => \_gnd_net_\
        );

    \cntr_RNIB8QE_2_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1762\,
            in1 => \N__1736\,
            in2 => \N__1670\,
            in3 => \N__1711\,
            lcout => un2_cntr_c4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_0_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2032\,
            lcout => \clk_divZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PORT_r_RNO_2_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1660\,
            in2 => \_gnd_net_\,
            in3 => \N__1624\,
            lcout => un1_cntr_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PORT_r_RNO_0_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001001"
        )
    port map (
            in0 => \N__1600\,
            in1 => \N__1576\,
            in2 => \N__1561\,
            in3 => \N__1533\,
            lcout => \PORT_r3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_11_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2095\,
            lcout => clk_div_i_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2187\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_1_cry_1_c_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2052\,
            in2 => \N__2035\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => clk_div_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_2_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2004\,
            in2 => \_gnd_net_\,
            in3 => \N__1990\,
            lcout => \clk_divZ0Z_2\,
            ltout => OPEN,
            carryin => clk_div_1_cry_1,
            carryout => clk_div_1_cry_2,
            clk => \N__2185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_3_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1986\,
            in2 => \_gnd_net_\,
            in3 => \N__1972\,
            lcout => \clk_divZ0Z_3\,
            ltout => OPEN,
            carryin => clk_div_1_cry_2,
            carryout => clk_div_1_cry_3,
            clk => \N__2185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_4_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1968\,
            in2 => \_gnd_net_\,
            in3 => \N__1954\,
            lcout => \clk_divZ0Z_4\,
            ltout => OPEN,
            carryin => clk_div_1_cry_3,
            carryout => clk_div_1_cry_4,
            clk => \N__2185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_5_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1950\,
            in2 => \_gnd_net_\,
            in3 => \N__1936\,
            lcout => \clk_divZ0Z_5\,
            ltout => OPEN,
            carryin => clk_div_1_cry_4,
            carryout => clk_div_1_cry_5,
            clk => \N__2185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_6_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1932\,
            in2 => \_gnd_net_\,
            in3 => \N__1918\,
            lcout => \clk_divZ0Z_6\,
            ltout => OPEN,
            carryin => clk_div_1_cry_5,
            carryout => clk_div_1_cry_6,
            clk => \N__2185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_7_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1914\,
            in2 => \_gnd_net_\,
            in3 => \N__1900\,
            lcout => \clk_divZ0Z_7\,
            ltout => OPEN,
            carryin => clk_div_1_cry_6,
            carryout => clk_div_1_cry_7,
            clk => \N__2185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_8_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2244\,
            in2 => \_gnd_net_\,
            in3 => \N__2230\,
            lcout => \clk_divZ0Z_8\,
            ltout => OPEN,
            carryin => clk_div_1_cry_7,
            carryout => clk_div_1_cry_8,
            clk => \N__2185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_9_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2226\,
            in2 => \_gnd_net_\,
            in3 => \N__2212\,
            lcout => \clk_divZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => clk_div_1_cry_9,
            clk => \N__2188\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_10_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2206\,
            in2 => \_gnd_net_\,
            in3 => \N__2209\,
            lcout => \clk_divZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2188\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \shift_ret_1_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__2519\,
            in1 => \_gnd_net_\,
            in2 => \N__2632\,
            in3 => \N__2573\,
            lcout => level_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \shift_0_2_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2627\,
            lcout => \shift_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \shift_0_1_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2518\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \shift_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2309\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \shift_ret_1_RNI69IQ_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__2574\,
            in1 => \N__2520\,
            in2 => \N__2592\,
            in3 => \N__2631\,
            lcout => \shift_ret_1_RNI69IQZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \up_2_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__2541\,
            in1 => \N__2148\,
            in2 => \_gnd_net_\,
            in3 => \N__2126\,
            lcout => \upZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2330\,
            ce => \N__2110\,
            sr => \_gnd_net_\
        );

    \up_1_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__2125\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2540\,
            lcout => \upZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2330\,
            ce => \N__2110\,
            sr => \_gnd_net_\
        );

    \up_e_0_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100011011001100"
        )
    port map (
            in0 => \N__2626\,
            in1 => \N__2539\,
            in2 => \N__2593\,
            in3 => \N__2575\,
            lcout => \upZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2325\,
            ce => \N__2521\,
            sr => \_gnd_net_\
        );

    \down_1_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2491\,
            in2 => \_gnd_net_\,
            in3 => \N__2361\,
            lcout => \downZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2334\,
            ce => \N__2455\,
            sr => \_gnd_net_\
        );

    \down_2_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__2466\,
            in1 => \N__2492\,
            in2 => \_gnd_net_\,
            in3 => \N__2362\,
            lcout => \downZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2334\,
            ce => \N__2455\,
            sr => \_gnd_net_\
        );

    \shift2_0_2_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2401\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \shift2_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \shift2_ret_1_RNITCI51_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__2439\,
            in1 => \N__2405\,
            in2 => \N__2428\,
            in3 => \N__2262\,
            lcout => \shift2_ret_1_RNITCIZ0Z51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \shift2_ret_1_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__2261\,
            in1 => \_gnd_net_\,
            in2 => \N__2409\,
            in3 => \N__2423\,
            lcout => level2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \shift2_0_1_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__2260\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \shift2_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2326\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \down_e_0_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011010011110000"
        )
    port map (
            in0 => \N__2440\,
            in1 => \N__2427\,
            in2 => \N__2369\,
            in3 => \N__2410\,
            lcout => \downZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2335\,
            ce => \N__2269\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
