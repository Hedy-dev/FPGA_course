// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jul 13 2021 15:22:48

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    LED5,
    LED1,
    LED6,
    LED4,
    LED2,
    LED0,
    CLK,
    LED7,
    LED3);

    output LED5;
    output LED1;
    output LED6;
    output LED4;
    output LED2;
    output LED0;
    input CLK;
    output LED7;
    output LED3;

    wire N__2484;
    wire N__2483;
    wire N__2482;
    wire N__2473;
    wire N__2472;
    wire N__2471;
    wire N__2464;
    wire N__2463;
    wire N__2462;
    wire N__2455;
    wire N__2454;
    wire N__2453;
    wire N__2446;
    wire N__2445;
    wire N__2444;
    wire N__2437;
    wire N__2436;
    wire N__2435;
    wire N__2428;
    wire N__2427;
    wire N__2426;
    wire N__2419;
    wire N__2418;
    wire N__2417;
    wire N__2410;
    wire N__2409;
    wire N__2408;
    wire N__2391;
    wire N__2390;
    wire N__2387;
    wire N__2384;
    wire N__2381;
    wire N__2376;
    wire N__2373;
    wire N__2372;
    wire N__2369;
    wire N__2366;
    wire N__2363;
    wire N__2358;
    wire N__2355;
    wire N__2354;
    wire N__2351;
    wire N__2348;
    wire N__2345;
    wire N__2340;
    wire N__2337;
    wire N__2336;
    wire N__2333;
    wire N__2330;
    wire N__2327;
    wire N__2322;
    wire N__2319;
    wire N__2318;
    wire N__2315;
    wire N__2312;
    wire N__2309;
    wire N__2304;
    wire N__2301;
    wire N__2300;
    wire N__2297;
    wire N__2294;
    wire N__2291;
    wire N__2286;
    wire N__2283;
    wire N__2280;
    wire N__2279;
    wire N__2276;
    wire N__2273;
    wire N__2268;
    wire N__2267;
    wire N__2266;
    wire N__2265;
    wire N__2264;
    wire N__2263;
    wire N__2262;
    wire N__2261;
    wire N__2244;
    wire N__2241;
    wire N__2238;
    wire N__2235;
    wire N__2234;
    wire N__2231;
    wire N__2228;
    wire N__2225;
    wire N__2220;
    wire N__2217;
    wire N__2216;
    wire N__2213;
    wire N__2210;
    wire N__2207;
    wire N__2202;
    wire N__2199;
    wire N__2198;
    wire N__2195;
    wire N__2192;
    wire N__2189;
    wire N__2184;
    wire N__2181;
    wire N__2180;
    wire N__2177;
    wire N__2174;
    wire N__2171;
    wire N__2166;
    wire N__2163;
    wire N__2162;
    wire N__2159;
    wire N__2156;
    wire N__2153;
    wire N__2148;
    wire N__2145;
    wire N__2144;
    wire N__2141;
    wire N__2138;
    wire N__2135;
    wire N__2130;
    wire N__2127;
    wire N__2126;
    wire N__2123;
    wire N__2120;
    wire N__2117;
    wire N__2112;
    wire N__2109;
    wire N__2108;
    wire N__2105;
    wire N__2102;
    wire N__2099;
    wire N__2094;
    wire N__2091;
    wire N__2090;
    wire N__2089;
    wire N__2086;
    wire N__2081;
    wire N__2076;
    wire N__2075;
    wire N__2072;
    wire N__2069;
    wire N__2064;
    wire N__2063;
    wire N__2062;
    wire N__2061;
    wire N__2060;
    wire N__2059;
    wire N__2058;
    wire N__2057;
    wire N__2054;
    wire N__2047;
    wire N__2042;
    wire N__2037;
    wire N__2028;
    wire N__2027;
    wire N__2024;
    wire N__2023;
    wire N__2022;
    wire N__2019;
    wire N__2016;
    wire N__2011;
    wire N__2004;
    wire N__2001;
    wire N__1998;
    wire N__1997;
    wire N__1996;
    wire N__1989;
    wire N__1988;
    wire N__1985;
    wire N__1982;
    wire N__1977;
    wire N__1976;
    wire N__1973;
    wire N__1970;
    wire N__1967;
    wire N__1966;
    wire N__1963;
    wire N__1960;
    wire N__1957;
    wire N__1954;
    wire N__1947;
    wire N__1946;
    wire N__1941;
    wire N__1938;
    wire N__1935;
    wire N__1932;
    wire N__1931;
    wire N__1930;
    wire N__1927;
    wire N__1926;
    wire N__1923;
    wire N__1922;
    wire N__1919;
    wire N__1916;
    wire N__1913;
    wire N__1908;
    wire N__1899;
    wire N__1896;
    wire N__1893;
    wire N__1890;
    wire N__1887;
    wire N__1884;
    wire N__1881;
    wire N__1880;
    wire N__1879;
    wire N__1876;
    wire N__1875;
    wire N__1872;
    wire N__1869;
    wire N__1866;
    wire N__1863;
    wire N__1860;
    wire N__1857;
    wire N__1854;
    wire N__1845;
    wire N__1842;
    wire N__1839;
    wire N__1836;
    wire N__1833;
    wire N__1832;
    wire N__1829;
    wire N__1828;
    wire N__1825;
    wire N__1822;
    wire N__1819;
    wire N__1816;
    wire N__1809;
    wire N__1808;
    wire N__1807;
    wire N__1806;
    wire N__1805;
    wire N__1804;
    wire N__1803;
    wire N__1802;
    wire N__1797;
    wire N__1794;
    wire N__1783;
    wire N__1776;
    wire N__1773;
    wire N__1770;
    wire N__1767;
    wire N__1766;
    wire N__1765;
    wire N__1764;
    wire N__1763;
    wire N__1762;
    wire N__1761;
    wire N__1758;
    wire N__1745;
    wire N__1740;
    wire N__1737;
    wire N__1736;
    wire N__1733;
    wire N__1730;
    wire N__1729;
    wire N__1726;
    wire N__1723;
    wire N__1720;
    wire N__1715;
    wire N__1710;
    wire N__1709;
    wire N__1706;
    wire N__1703;
    wire N__1700;
    wire N__1697;
    wire N__1694;
    wire N__1689;
    wire N__1688;
    wire N__1685;
    wire N__1684;
    wire N__1681;
    wire N__1678;
    wire N__1675;
    wire N__1668;
    wire N__1665;
    wire N__1664;
    wire N__1663;
    wire N__1662;
    wire N__1659;
    wire N__1656;
    wire N__1651;
    wire N__1648;
    wire N__1645;
    wire N__1638;
    wire N__1637;
    wire N__1634;
    wire N__1631;
    wire N__1628;
    wire N__1623;
    wire N__1620;
    wire N__1619;
    wire N__1616;
    wire N__1613;
    wire N__1610;
    wire N__1605;
    wire N__1602;
    wire N__1599;
    wire N__1596;
    wire N__1595;
    wire N__1594;
    wire N__1593;
    wire N__1592;
    wire N__1589;
    wire N__1588;
    wire N__1587;
    wire N__1584;
    wire N__1579;
    wire N__1574;
    wire N__1569;
    wire N__1560;
    wire N__1557;
    wire N__1556;
    wire N__1553;
    wire N__1550;
    wire N__1545;
    wire N__1544;
    wire N__1543;
    wire N__1542;
    wire N__1541;
    wire N__1538;
    wire N__1535;
    wire N__1532;
    wire N__1527;
    wire N__1518;
    wire N__1515;
    wire N__1514;
    wire N__1511;
    wire N__1510;
    wire N__1509;
    wire N__1508;
    wire N__1507;
    wire N__1506;
    wire N__1505;
    wire N__1502;
    wire N__1499;
    wire N__1494;
    wire N__1489;
    wire N__1484;
    wire N__1473;
    wire N__1472;
    wire N__1471;
    wire N__1470;
    wire N__1469;
    wire N__1466;
    wire N__1463;
    wire N__1458;
    wire N__1455;
    wire N__1446;
    wire N__1443;
    wire N__1442;
    wire N__1441;
    wire N__1440;
    wire N__1437;
    wire N__1434;
    wire N__1427;
    wire N__1422;
    wire N__1421;
    wire N__1420;
    wire N__1419;
    wire N__1410;
    wire N__1407;
    wire N__1406;
    wire N__1405;
    wire N__1402;
    wire N__1399;
    wire N__1396;
    wire N__1389;
    wire N__1386;
    wire N__1383;
    wire N__1382;
    wire N__1377;
    wire N__1374;
    wire N__1371;
    wire N__1370;
    wire N__1369;
    wire N__1368;
    wire N__1367;
    wire N__1364;
    wire N__1361;
    wire N__1356;
    wire N__1353;
    wire N__1344;
    wire N__1341;
    wire N__1338;
    wire N__1335;
    wire N__1332;
    wire N__1329;
    wire N__1326;
    wire N__1323;
    wire N__1320;
    wire N__1317;
    wire N__1316;
    wire N__1313;
    wire N__1310;
    wire N__1309;
    wire N__1306;
    wire N__1303;
    wire N__1300;
    wire N__1293;
    wire N__1290;
    wire N__1287;
    wire N__1284;
    wire N__1281;
    wire N__1280;
    wire N__1277;
    wire N__1274;
    wire N__1273;
    wire N__1270;
    wire N__1267;
    wire N__1264;
    wire N__1261;
    wire N__1256;
    wire N__1251;
    wire N__1248;
    wire N__1245;
    wire N__1242;
    wire N__1241;
    wire N__1238;
    wire N__1235;
    wire N__1234;
    wire N__1231;
    wire N__1228;
    wire N__1225;
    wire N__1218;
    wire N__1215;
    wire N__1212;
    wire N__1209;
    wire N__1206;
    wire N__1205;
    wire N__1202;
    wire N__1199;
    wire N__1198;
    wire N__1195;
    wire N__1192;
    wire N__1189;
    wire N__1182;
    wire N__1179;
    wire N__1176;
    wire N__1175;
    wire N__1172;
    wire N__1169;
    wire N__1168;
    wire N__1165;
    wire N__1162;
    wire N__1159;
    wire N__1152;
    wire N__1149;
    wire N__1146;
    wire N__1143;
    wire N__1140;
    wire N__1137;
    wire N__1134;
    wire N__1131;
    wire N__1130;
    wire N__1125;
    wire N__1122;
    wire N__1119;
    wire GNDG0;
    wire VCCG0;
    wire BIT_47_0_a3_0_1_6_cascade_;
    wire N_17_cascade_;
    wire N_22_cascade_;
    wire BIT_47_0_a3_0_1_6;
    wire N_31;
    wire BIT_47_0;
    wire LED0_c;
    wire clk_div_RNIICCP5Z0Z_19_cascade_;
    wire N_12_i;
    wire LED2_c;
    wire N_14_i;
    wire LED3_c;
    wire N_6_i;
    wire LED4_c;
    wire N_8_i;
    wire LED5_c;
    wire bfn_1_8_0_;
    wire clk_div_2_cry_1;
    wire clk_div_2_cry_2;
    wire clk_div_2_cry_3;
    wire clk_div_2_cry_4;
    wire clk_div_2_cry_5;
    wire clk_div_2_cry_6;
    wire clk_div_2_cry_7;
    wire clk_div_2_cry_8;
    wire bfn_1_9_0_;
    wire clk_div_2_cry_9;
    wire clk_div_2_cry_10;
    wire clk_div_2_cry_11;
    wire clk_div_2_cry_12;
    wire clk_div_2_cry_13;
    wire clk_div_2_cry_14;
    wire clk_div_2_cry_15;
    wire clk_div_2_cry_16;
    wire bfn_1_10_0_;
    wire clk_div_2_cry_17;
    wire clk_div_2_cry_18;
    wire BIT_47_i_o3_0_0_4_cascade_;
    wire N_27;
    wire N_45;
    wire N_17;
    wire N_45_cascade_;
    wire N_30;
    wire bfn_2_6_0_;
    wire cntrZ0Z_1;
    wire cntr_cry_0;
    wire cntr_cry_1;
    wire cntr_cry_2;
    wire cntr_cry_3;
    wire cntr_cry_4;
    wire cntr_cry_5;
    wire cntrZ0Z_6;
    wire N_23;
    wire cntrZ0Z_2;
    wire N_21_cascade_;
    wire cntrZ0Z_5;
    wire cntrZ0Z_0;
    wire clk_div_i_19;
    wire cntrZ0Z_3;
    wire N_22;
    wire N_21;
    wire N_19;
    wire LED1_c;
    wire N_38;
    wire BIT_47_1;
    wire cntrZ0Z_4;
    wire g0_0;
    wire g0_4;
    wire clk_div_RNIK8D95Z0Z_19;
    wire cntr_RNIVLLQ5Z0Z_4_cascade_;
    wire BIT_47_6;
    wire LED6_c;
    wire clk_div_RNIICCP5Z0Z_19;
    wire BIT_47_7;
    wire cntr_RNIVLLQ5Z0Z_4;
    wire LED7_c;
    wire clk_div_RNI0HSQ5Z0Z_19;
    wire clk_divZ0Z_1;
    wire clk_divZ0Z_0;
    wire bfn_2_9_0_;
    wire clk_divZ0Z_2;
    wire clk_div_1_cry_1;
    wire clk_divZ0Z_3;
    wire clk_div_1_cry_2;
    wire clk_divZ0Z_4;
    wire clk_div_1_cry_3;
    wire clk_divZ0Z_5;
    wire clk_div_1_cry_4;
    wire clk_divZ0Z_6;
    wire clk_div_1_cry_5;
    wire clk_divZ0Z_7;
    wire clk_div_1_cry_6;
    wire clk_divZ0Z_8;
    wire clk_div_1_cry_7;
    wire clk_div_1_cry_8;
    wire clk_divZ0Z_9;
    wire bfn_2_10_0_;
    wire clk_divZ0Z_10;
    wire clk_div_1_cry_9;
    wire clk_divZ0Z_11;
    wire clk_div_1_cry_10;
    wire clk_divZ0Z_12;
    wire clk_div_1_cry_11;
    wire clk_divZ0Z_13;
    wire clk_div_1_cry_12;
    wire clk_divZ0Z_14;
    wire clk_div_1_cry_13;
    wire clk_divZ0Z_15;
    wire clk_div_1_cry_14;
    wire clk_divZ0Z_16;
    wire clk_div_1_cry_15;
    wire clk_div_1_cry_16;
    wire clk_divZ0Z_17;
    wire bfn_2_11_0_;
    wire clk_div_1_cry_17;
    wire clk_divZ0Z_18;
    wire CLK_0_c_g;
    wire _gnd_net_;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__2482),
            .GLOBALBUFFEROUTPUT(CLK_0_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__2484),
            .DIN(N__2483),
            .DOUT(N__2482),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__2484),
            .PADOUT(N__2483),
            .PADIN(N__2482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED4_obuf_iopad (
            .OE(N__2473),
            .DIN(N__2472),
            .DOUT(N__2471),
            .PACKAGEPIN(LED4));
    defparam LED4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED4_obuf_preio (
            .PADOEN(N__2473),
            .PADOUT(N__2472),
            .PADIN(N__2471),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1212),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED2_obuf_iopad (
            .OE(N__2464),
            .DIN(N__2463),
            .DOUT(N__2462),
            .PACKAGEPIN(LED2));
    defparam LED2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED2_obuf_preio (
            .PADOEN(N__2464),
            .PADOUT(N__2463),
            .PADIN(N__2462),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1284),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED0_obuf_iopad (
            .OE(N__2455),
            .DIN(N__2454),
            .DOUT(N__2453),
            .PACKAGEPIN(LED0));
    defparam LED0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED0_obuf_preio (
            .PADOEN(N__2455),
            .PADOUT(N__2454),
            .PADIN(N__2453),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1326),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED6_obuf_iopad (
            .OE(N__2446),
            .DIN(N__2445),
            .DOUT(N__2444),
            .PACKAGEPIN(LED6));
    defparam LED6_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED6_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED6_obuf_preio (
            .PADOEN(N__2446),
            .PADOUT(N__2445),
            .PADIN(N__2444),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1836),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED3_obuf_iopad (
            .OE(N__2437),
            .DIN(N__2436),
            .DOUT(N__2435),
            .PACKAGEPIN(LED3));
    defparam LED3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED3_obuf_preio (
            .PADOEN(N__2437),
            .PADOUT(N__2436),
            .PADIN(N__2435),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1245),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED7_obuf_iopad (
            .OE(N__2428),
            .DIN(N__2427),
            .DOUT(N__2426),
            .PACKAGEPIN(LED7));
    defparam LED7_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED7_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED7_obuf_preio (
            .PADOEN(N__2428),
            .PADOUT(N__2427),
            .PADIN(N__2426),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1740),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED1_obuf_iopad (
            .OE(N__2419),
            .DIN(N__2418),
            .DOUT(N__2417),
            .PACKAGEPIN(LED1));
    defparam LED1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED1_obuf_preio (
            .PADOEN(N__2419),
            .PADOUT(N__2418),
            .PADIN(N__2417),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1977),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED5_obuf_iopad (
            .OE(N__2410),
            .DIN(N__2409),
            .DOUT(N__2408),
            .PACKAGEPIN(LED5));
    defparam LED5_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED5_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED5_obuf_preio (
            .PADOEN(N__2410),
            .PADOUT(N__2409),
            .PADIN(N__2408),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1176),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__523 (
            .O(N__2391),
            .I(N__2387));
    InMux I__522 (
            .O(N__2390),
            .I(N__2384));
    InMux I__521 (
            .O(N__2387),
            .I(N__2381));
    LocalMux I__520 (
            .O(N__2384),
            .I(clk_divZ0Z_12));
    LocalMux I__519 (
            .O(N__2381),
            .I(clk_divZ0Z_12));
    InMux I__518 (
            .O(N__2376),
            .I(clk_div_1_cry_11));
    CascadeMux I__517 (
            .O(N__2373),
            .I(N__2369));
    InMux I__516 (
            .O(N__2372),
            .I(N__2366));
    InMux I__515 (
            .O(N__2369),
            .I(N__2363));
    LocalMux I__514 (
            .O(N__2366),
            .I(clk_divZ0Z_13));
    LocalMux I__513 (
            .O(N__2363),
            .I(clk_divZ0Z_13));
    InMux I__512 (
            .O(N__2358),
            .I(clk_div_1_cry_12));
    CascadeMux I__511 (
            .O(N__2355),
            .I(N__2351));
    InMux I__510 (
            .O(N__2354),
            .I(N__2348));
    InMux I__509 (
            .O(N__2351),
            .I(N__2345));
    LocalMux I__508 (
            .O(N__2348),
            .I(clk_divZ0Z_14));
    LocalMux I__507 (
            .O(N__2345),
            .I(clk_divZ0Z_14));
    InMux I__506 (
            .O(N__2340),
            .I(clk_div_1_cry_13));
    CascadeMux I__505 (
            .O(N__2337),
            .I(N__2333));
    InMux I__504 (
            .O(N__2336),
            .I(N__2330));
    InMux I__503 (
            .O(N__2333),
            .I(N__2327));
    LocalMux I__502 (
            .O(N__2330),
            .I(clk_divZ0Z_15));
    LocalMux I__501 (
            .O(N__2327),
            .I(clk_divZ0Z_15));
    InMux I__500 (
            .O(N__2322),
            .I(clk_div_1_cry_14));
    CascadeMux I__499 (
            .O(N__2319),
            .I(N__2315));
    InMux I__498 (
            .O(N__2318),
            .I(N__2312));
    InMux I__497 (
            .O(N__2315),
            .I(N__2309));
    LocalMux I__496 (
            .O(N__2312),
            .I(clk_divZ0Z_16));
    LocalMux I__495 (
            .O(N__2309),
            .I(clk_divZ0Z_16));
    InMux I__494 (
            .O(N__2304),
            .I(clk_div_1_cry_15));
    CascadeMux I__493 (
            .O(N__2301),
            .I(N__2297));
    InMux I__492 (
            .O(N__2300),
            .I(N__2294));
    InMux I__491 (
            .O(N__2297),
            .I(N__2291));
    LocalMux I__490 (
            .O(N__2294),
            .I(clk_divZ0Z_17));
    LocalMux I__489 (
            .O(N__2291),
            .I(clk_divZ0Z_17));
    InMux I__488 (
            .O(N__2286),
            .I(bfn_2_11_0_));
    InMux I__487 (
            .O(N__2283),
            .I(clk_div_1_cry_17));
    InMux I__486 (
            .O(N__2280),
            .I(N__2276));
    InMux I__485 (
            .O(N__2279),
            .I(N__2273));
    LocalMux I__484 (
            .O(N__2276),
            .I(clk_divZ0Z_18));
    LocalMux I__483 (
            .O(N__2273),
            .I(clk_divZ0Z_18));
    ClkMux I__482 (
            .O(N__2268),
            .I(N__2244));
    ClkMux I__481 (
            .O(N__2267),
            .I(N__2244));
    ClkMux I__480 (
            .O(N__2266),
            .I(N__2244));
    ClkMux I__479 (
            .O(N__2265),
            .I(N__2244));
    ClkMux I__478 (
            .O(N__2264),
            .I(N__2244));
    ClkMux I__477 (
            .O(N__2263),
            .I(N__2244));
    ClkMux I__476 (
            .O(N__2262),
            .I(N__2244));
    ClkMux I__475 (
            .O(N__2261),
            .I(N__2244));
    GlobalMux I__474 (
            .O(N__2244),
            .I(N__2241));
    gio2CtrlBuf I__473 (
            .O(N__2241),
            .I(CLK_0_c_g));
    InMux I__472 (
            .O(N__2238),
            .I(clk_div_1_cry_2));
    CascadeMux I__471 (
            .O(N__2235),
            .I(N__2231));
    InMux I__470 (
            .O(N__2234),
            .I(N__2228));
    InMux I__469 (
            .O(N__2231),
            .I(N__2225));
    LocalMux I__468 (
            .O(N__2228),
            .I(clk_divZ0Z_4));
    LocalMux I__467 (
            .O(N__2225),
            .I(clk_divZ0Z_4));
    InMux I__466 (
            .O(N__2220),
            .I(clk_div_1_cry_3));
    CascadeMux I__465 (
            .O(N__2217),
            .I(N__2213));
    InMux I__464 (
            .O(N__2216),
            .I(N__2210));
    InMux I__463 (
            .O(N__2213),
            .I(N__2207));
    LocalMux I__462 (
            .O(N__2210),
            .I(clk_divZ0Z_5));
    LocalMux I__461 (
            .O(N__2207),
            .I(clk_divZ0Z_5));
    InMux I__460 (
            .O(N__2202),
            .I(clk_div_1_cry_4));
    CascadeMux I__459 (
            .O(N__2199),
            .I(N__2195));
    InMux I__458 (
            .O(N__2198),
            .I(N__2192));
    InMux I__457 (
            .O(N__2195),
            .I(N__2189));
    LocalMux I__456 (
            .O(N__2192),
            .I(clk_divZ0Z_6));
    LocalMux I__455 (
            .O(N__2189),
            .I(clk_divZ0Z_6));
    InMux I__454 (
            .O(N__2184),
            .I(clk_div_1_cry_5));
    CascadeMux I__453 (
            .O(N__2181),
            .I(N__2177));
    InMux I__452 (
            .O(N__2180),
            .I(N__2174));
    InMux I__451 (
            .O(N__2177),
            .I(N__2171));
    LocalMux I__450 (
            .O(N__2174),
            .I(clk_divZ0Z_7));
    LocalMux I__449 (
            .O(N__2171),
            .I(clk_divZ0Z_7));
    InMux I__448 (
            .O(N__2166),
            .I(clk_div_1_cry_6));
    CascadeMux I__447 (
            .O(N__2163),
            .I(N__2159));
    InMux I__446 (
            .O(N__2162),
            .I(N__2156));
    InMux I__445 (
            .O(N__2159),
            .I(N__2153));
    LocalMux I__444 (
            .O(N__2156),
            .I(clk_divZ0Z_8));
    LocalMux I__443 (
            .O(N__2153),
            .I(clk_divZ0Z_8));
    InMux I__442 (
            .O(N__2148),
            .I(clk_div_1_cry_7));
    CascadeMux I__441 (
            .O(N__2145),
            .I(N__2141));
    InMux I__440 (
            .O(N__2144),
            .I(N__2138));
    InMux I__439 (
            .O(N__2141),
            .I(N__2135));
    LocalMux I__438 (
            .O(N__2138),
            .I(clk_divZ0Z_9));
    LocalMux I__437 (
            .O(N__2135),
            .I(clk_divZ0Z_9));
    InMux I__436 (
            .O(N__2130),
            .I(bfn_2_10_0_));
    CascadeMux I__435 (
            .O(N__2127),
            .I(N__2123));
    InMux I__434 (
            .O(N__2126),
            .I(N__2120));
    InMux I__433 (
            .O(N__2123),
            .I(N__2117));
    LocalMux I__432 (
            .O(N__2120),
            .I(clk_divZ0Z_10));
    LocalMux I__431 (
            .O(N__2117),
            .I(clk_divZ0Z_10));
    InMux I__430 (
            .O(N__2112),
            .I(clk_div_1_cry_9));
    CascadeMux I__429 (
            .O(N__2109),
            .I(N__2105));
    InMux I__428 (
            .O(N__2108),
            .I(N__2102));
    InMux I__427 (
            .O(N__2105),
            .I(N__2099));
    LocalMux I__426 (
            .O(N__2102),
            .I(clk_divZ0Z_11));
    LocalMux I__425 (
            .O(N__2099),
            .I(clk_divZ0Z_11));
    InMux I__424 (
            .O(N__2094),
            .I(clk_div_1_cry_10));
    InMux I__423 (
            .O(N__2091),
            .I(N__2086));
    InMux I__422 (
            .O(N__2090),
            .I(N__2081));
    InMux I__421 (
            .O(N__2089),
            .I(N__2081));
    LocalMux I__420 (
            .O(N__2086),
            .I(N__2076));
    LocalMux I__419 (
            .O(N__2081),
            .I(N__2076));
    Span4Mux_h I__418 (
            .O(N__2076),
            .I(N__2072));
    InMux I__417 (
            .O(N__2075),
            .I(N__2069));
    Odrv4 I__416 (
            .O(N__2072),
            .I(clk_div_i_19));
    LocalMux I__415 (
            .O(N__2069),
            .I(clk_div_i_19));
    InMux I__414 (
            .O(N__2064),
            .I(N__2054));
    InMux I__413 (
            .O(N__2063),
            .I(N__2047));
    InMux I__412 (
            .O(N__2062),
            .I(N__2047));
    InMux I__411 (
            .O(N__2061),
            .I(N__2047));
    InMux I__410 (
            .O(N__2060),
            .I(N__2042));
    InMux I__409 (
            .O(N__2059),
            .I(N__2042));
    InMux I__408 (
            .O(N__2058),
            .I(N__2037));
    InMux I__407 (
            .O(N__2057),
            .I(N__2037));
    LocalMux I__406 (
            .O(N__2054),
            .I(cntrZ0Z_3));
    LocalMux I__405 (
            .O(N__2047),
            .I(cntrZ0Z_3));
    LocalMux I__404 (
            .O(N__2042),
            .I(cntrZ0Z_3));
    LocalMux I__403 (
            .O(N__2037),
            .I(cntrZ0Z_3));
    CascadeMux I__402 (
            .O(N__2028),
            .I(N__2024));
    InMux I__401 (
            .O(N__2027),
            .I(N__2019));
    InMux I__400 (
            .O(N__2024),
            .I(N__2016));
    InMux I__399 (
            .O(N__2023),
            .I(N__2011));
    InMux I__398 (
            .O(N__2022),
            .I(N__2011));
    LocalMux I__397 (
            .O(N__2019),
            .I(N_22));
    LocalMux I__396 (
            .O(N__2016),
            .I(N_22));
    LocalMux I__395 (
            .O(N__2011),
            .I(N_22));
    InMux I__394 (
            .O(N__2004),
            .I(N__2001));
    LocalMux I__393 (
            .O(N__2001),
            .I(N_21));
    InMux I__392 (
            .O(N__1998),
            .I(N__1989));
    InMux I__391 (
            .O(N__1997),
            .I(N__1989));
    InMux I__390 (
            .O(N__1996),
            .I(N__1989));
    LocalMux I__389 (
            .O(N__1989),
            .I(N__1985));
    InMux I__388 (
            .O(N__1988),
            .I(N__1982));
    Odrv4 I__387 (
            .O(N__1985),
            .I(N_19));
    LocalMux I__386 (
            .O(N__1982),
            .I(N_19));
    IoInMux I__385 (
            .O(N__1977),
            .I(N__1973));
    CascadeMux I__384 (
            .O(N__1976),
            .I(N__1970));
    LocalMux I__383 (
            .O(N__1973),
            .I(N__1967));
    InMux I__382 (
            .O(N__1970),
            .I(N__1963));
    Span4Mux_s0_h I__381 (
            .O(N__1967),
            .I(N__1960));
    InMux I__380 (
            .O(N__1966),
            .I(N__1957));
    LocalMux I__379 (
            .O(N__1963),
            .I(N__1954));
    Odrv4 I__378 (
            .O(N__1960),
            .I(LED1_c));
    LocalMux I__377 (
            .O(N__1957),
            .I(LED1_c));
    Odrv4 I__376 (
            .O(N__1954),
            .I(LED1_c));
    InMux I__375 (
            .O(N__1947),
            .I(N__1941));
    InMux I__374 (
            .O(N__1946),
            .I(N__1941));
    LocalMux I__373 (
            .O(N__1941),
            .I(N_38));
    InMux I__372 (
            .O(N__1938),
            .I(N__1935));
    LocalMux I__371 (
            .O(N__1935),
            .I(BIT_47_1));
    InMux I__370 (
            .O(N__1932),
            .I(N__1927));
    CascadeMux I__369 (
            .O(N__1931),
            .I(N__1923));
    InMux I__368 (
            .O(N__1930),
            .I(N__1919));
    LocalMux I__367 (
            .O(N__1927),
            .I(N__1916));
    InMux I__366 (
            .O(N__1926),
            .I(N__1913));
    InMux I__365 (
            .O(N__1923),
            .I(N__1908));
    InMux I__364 (
            .O(N__1922),
            .I(N__1908));
    LocalMux I__363 (
            .O(N__1919),
            .I(cntrZ0Z_4));
    Odrv4 I__362 (
            .O(N__1916),
            .I(cntrZ0Z_4));
    LocalMux I__361 (
            .O(N__1913),
            .I(cntrZ0Z_4));
    LocalMux I__360 (
            .O(N__1908),
            .I(cntrZ0Z_4));
    InMux I__359 (
            .O(N__1899),
            .I(N__1896));
    LocalMux I__358 (
            .O(N__1896),
            .I(N__1893));
    Odrv4 I__357 (
            .O(N__1893),
            .I(g0_0));
    CascadeMux I__356 (
            .O(N__1890),
            .I(N__1887));
    InMux I__355 (
            .O(N__1887),
            .I(N__1884));
    LocalMux I__354 (
            .O(N__1884),
            .I(g0_4));
    CascadeMux I__353 (
            .O(N__1881),
            .I(N__1876));
    InMux I__352 (
            .O(N__1880),
            .I(N__1872));
    InMux I__351 (
            .O(N__1879),
            .I(N__1869));
    InMux I__350 (
            .O(N__1876),
            .I(N__1866));
    InMux I__349 (
            .O(N__1875),
            .I(N__1863));
    LocalMux I__348 (
            .O(N__1872),
            .I(N__1860));
    LocalMux I__347 (
            .O(N__1869),
            .I(N__1857));
    LocalMux I__346 (
            .O(N__1866),
            .I(N__1854));
    LocalMux I__345 (
            .O(N__1863),
            .I(clk_div_RNIK8D95Z0Z_19));
    Odrv4 I__344 (
            .O(N__1860),
            .I(clk_div_RNIK8D95Z0Z_19));
    Odrv4 I__343 (
            .O(N__1857),
            .I(clk_div_RNIK8D95Z0Z_19));
    Odrv4 I__342 (
            .O(N__1854),
            .I(clk_div_RNIK8D95Z0Z_19));
    CascadeMux I__341 (
            .O(N__1845),
            .I(cntr_RNIVLLQ5Z0Z_4_cascade_));
    InMux I__340 (
            .O(N__1842),
            .I(N__1839));
    LocalMux I__339 (
            .O(N__1839),
            .I(BIT_47_6));
    IoInMux I__338 (
            .O(N__1836),
            .I(N__1833));
    LocalMux I__337 (
            .O(N__1833),
            .I(N__1829));
    InMux I__336 (
            .O(N__1832),
            .I(N__1825));
    Span4Mux_s3_v I__335 (
            .O(N__1829),
            .I(N__1822));
    InMux I__334 (
            .O(N__1828),
            .I(N__1819));
    LocalMux I__333 (
            .O(N__1825),
            .I(N__1816));
    Odrv4 I__332 (
            .O(N__1822),
            .I(LED6_c));
    LocalMux I__331 (
            .O(N__1819),
            .I(LED6_c));
    Odrv4 I__330 (
            .O(N__1816),
            .I(LED6_c));
    InMux I__329 (
            .O(N__1809),
            .I(N__1797));
    InMux I__328 (
            .O(N__1808),
            .I(N__1797));
    CEMux I__327 (
            .O(N__1807),
            .I(N__1794));
    InMux I__326 (
            .O(N__1806),
            .I(N__1783));
    InMux I__325 (
            .O(N__1805),
            .I(N__1783));
    InMux I__324 (
            .O(N__1804),
            .I(N__1783));
    InMux I__323 (
            .O(N__1803),
            .I(N__1783));
    InMux I__322 (
            .O(N__1802),
            .I(N__1783));
    LocalMux I__321 (
            .O(N__1797),
            .I(clk_div_RNIICCP5Z0Z_19));
    LocalMux I__320 (
            .O(N__1794),
            .I(clk_div_RNIICCP5Z0Z_19));
    LocalMux I__319 (
            .O(N__1783),
            .I(clk_div_RNIICCP5Z0Z_19));
    CascadeMux I__318 (
            .O(N__1776),
            .I(N__1773));
    InMux I__317 (
            .O(N__1773),
            .I(N__1770));
    LocalMux I__316 (
            .O(N__1770),
            .I(BIT_47_7));
    InMux I__315 (
            .O(N__1767),
            .I(N__1758));
    InMux I__314 (
            .O(N__1766),
            .I(N__1745));
    InMux I__313 (
            .O(N__1765),
            .I(N__1745));
    InMux I__312 (
            .O(N__1764),
            .I(N__1745));
    InMux I__311 (
            .O(N__1763),
            .I(N__1745));
    InMux I__310 (
            .O(N__1762),
            .I(N__1745));
    InMux I__309 (
            .O(N__1761),
            .I(N__1745));
    LocalMux I__308 (
            .O(N__1758),
            .I(cntr_RNIVLLQ5Z0Z_4));
    LocalMux I__307 (
            .O(N__1745),
            .I(cntr_RNIVLLQ5Z0Z_4));
    IoInMux I__306 (
            .O(N__1740),
            .I(N__1737));
    LocalMux I__305 (
            .O(N__1737),
            .I(N__1733));
    CascadeMux I__304 (
            .O(N__1736),
            .I(N__1730));
    IoSpan4Mux I__303 (
            .O(N__1733),
            .I(N__1726));
    InMux I__302 (
            .O(N__1730),
            .I(N__1723));
    InMux I__301 (
            .O(N__1729),
            .I(N__1720));
    Span4Mux_s1_h I__300 (
            .O(N__1726),
            .I(N__1715));
    LocalMux I__299 (
            .O(N__1723),
            .I(N__1715));
    LocalMux I__298 (
            .O(N__1720),
            .I(LED7_c));
    Odrv4 I__297 (
            .O(N__1715),
            .I(LED7_c));
    SRMux I__296 (
            .O(N__1710),
            .I(N__1706));
    SRMux I__295 (
            .O(N__1709),
            .I(N__1703));
    LocalMux I__294 (
            .O(N__1706),
            .I(N__1700));
    LocalMux I__293 (
            .O(N__1703),
            .I(N__1697));
    Span4Mux_s2_h I__292 (
            .O(N__1700),
            .I(N__1694));
    Odrv4 I__291 (
            .O(N__1697),
            .I(clk_div_RNI0HSQ5Z0Z_19));
    Odrv4 I__290 (
            .O(N__1694),
            .I(clk_div_RNI0HSQ5Z0Z_19));
    InMux I__289 (
            .O(N__1689),
            .I(N__1685));
    InMux I__288 (
            .O(N__1688),
            .I(N__1681));
    LocalMux I__287 (
            .O(N__1685),
            .I(N__1678));
    InMux I__286 (
            .O(N__1684),
            .I(N__1675));
    LocalMux I__285 (
            .O(N__1681),
            .I(clk_divZ0Z_1));
    Odrv4 I__284 (
            .O(N__1678),
            .I(clk_divZ0Z_1));
    LocalMux I__283 (
            .O(N__1675),
            .I(clk_divZ0Z_1));
    CascadeMux I__282 (
            .O(N__1668),
            .I(N__1665));
    InMux I__281 (
            .O(N__1665),
            .I(N__1659));
    CascadeMux I__280 (
            .O(N__1664),
            .I(N__1656));
    InMux I__279 (
            .O(N__1663),
            .I(N__1651));
    InMux I__278 (
            .O(N__1662),
            .I(N__1651));
    LocalMux I__277 (
            .O(N__1659),
            .I(N__1648));
    InMux I__276 (
            .O(N__1656),
            .I(N__1645));
    LocalMux I__275 (
            .O(N__1651),
            .I(clk_divZ0Z_0));
    Odrv4 I__274 (
            .O(N__1648),
            .I(clk_divZ0Z_0));
    LocalMux I__273 (
            .O(N__1645),
            .I(clk_divZ0Z_0));
    CascadeMux I__272 (
            .O(N__1638),
            .I(N__1634));
    InMux I__271 (
            .O(N__1637),
            .I(N__1631));
    InMux I__270 (
            .O(N__1634),
            .I(N__1628));
    LocalMux I__269 (
            .O(N__1631),
            .I(clk_divZ0Z_2));
    LocalMux I__268 (
            .O(N__1628),
            .I(clk_divZ0Z_2));
    InMux I__267 (
            .O(N__1623),
            .I(clk_div_1_cry_1));
    CascadeMux I__266 (
            .O(N__1620),
            .I(N__1616));
    InMux I__265 (
            .O(N__1619),
            .I(N__1613));
    InMux I__264 (
            .O(N__1616),
            .I(N__1610));
    LocalMux I__263 (
            .O(N__1613),
            .I(clk_divZ0Z_3));
    LocalMux I__262 (
            .O(N__1610),
            .I(clk_divZ0Z_3));
    InMux I__261 (
            .O(N__1605),
            .I(cntr_cry_3));
    InMux I__260 (
            .O(N__1602),
            .I(cntr_cry_4));
    InMux I__259 (
            .O(N__1599),
            .I(cntr_cry_5));
    CascadeMux I__258 (
            .O(N__1596),
            .I(N__1589));
    InMux I__257 (
            .O(N__1595),
            .I(N__1584));
    InMux I__256 (
            .O(N__1594),
            .I(N__1579));
    InMux I__255 (
            .O(N__1593),
            .I(N__1579));
    InMux I__254 (
            .O(N__1592),
            .I(N__1574));
    InMux I__253 (
            .O(N__1589),
            .I(N__1574));
    InMux I__252 (
            .O(N__1588),
            .I(N__1569));
    InMux I__251 (
            .O(N__1587),
            .I(N__1569));
    LocalMux I__250 (
            .O(N__1584),
            .I(cntrZ0Z_6));
    LocalMux I__249 (
            .O(N__1579),
            .I(cntrZ0Z_6));
    LocalMux I__248 (
            .O(N__1574),
            .I(cntrZ0Z_6));
    LocalMux I__247 (
            .O(N__1569),
            .I(cntrZ0Z_6));
    InMux I__246 (
            .O(N__1560),
            .I(N__1557));
    LocalMux I__245 (
            .O(N__1557),
            .I(N__1553));
    InMux I__244 (
            .O(N__1556),
            .I(N__1550));
    Odrv4 I__243 (
            .O(N__1553),
            .I(N_23));
    LocalMux I__242 (
            .O(N__1550),
            .I(N_23));
    InMux I__241 (
            .O(N__1545),
            .I(N__1538));
    InMux I__240 (
            .O(N__1544),
            .I(N__1535));
    InMux I__239 (
            .O(N__1543),
            .I(N__1532));
    InMux I__238 (
            .O(N__1542),
            .I(N__1527));
    InMux I__237 (
            .O(N__1541),
            .I(N__1527));
    LocalMux I__236 (
            .O(N__1538),
            .I(cntrZ0Z_2));
    LocalMux I__235 (
            .O(N__1535),
            .I(cntrZ0Z_2));
    LocalMux I__234 (
            .O(N__1532),
            .I(cntrZ0Z_2));
    LocalMux I__233 (
            .O(N__1527),
            .I(cntrZ0Z_2));
    CascadeMux I__232 (
            .O(N__1518),
            .I(N_21_cascade_));
    CascadeMux I__231 (
            .O(N__1515),
            .I(N__1511));
    InMux I__230 (
            .O(N__1514),
            .I(N__1502));
    InMux I__229 (
            .O(N__1511),
            .I(N__1499));
    InMux I__228 (
            .O(N__1510),
            .I(N__1494));
    InMux I__227 (
            .O(N__1509),
            .I(N__1494));
    InMux I__226 (
            .O(N__1508),
            .I(N__1489));
    InMux I__225 (
            .O(N__1507),
            .I(N__1489));
    InMux I__224 (
            .O(N__1506),
            .I(N__1484));
    InMux I__223 (
            .O(N__1505),
            .I(N__1484));
    LocalMux I__222 (
            .O(N__1502),
            .I(cntrZ0Z_5));
    LocalMux I__221 (
            .O(N__1499),
            .I(cntrZ0Z_5));
    LocalMux I__220 (
            .O(N__1494),
            .I(cntrZ0Z_5));
    LocalMux I__219 (
            .O(N__1489),
            .I(cntrZ0Z_5));
    LocalMux I__218 (
            .O(N__1484),
            .I(cntrZ0Z_5));
    InMux I__217 (
            .O(N__1473),
            .I(N__1466));
    InMux I__216 (
            .O(N__1472),
            .I(N__1463));
    InMux I__215 (
            .O(N__1471),
            .I(N__1458));
    InMux I__214 (
            .O(N__1470),
            .I(N__1458));
    InMux I__213 (
            .O(N__1469),
            .I(N__1455));
    LocalMux I__212 (
            .O(N__1466),
            .I(cntrZ0Z_0));
    LocalMux I__211 (
            .O(N__1463),
            .I(cntrZ0Z_0));
    LocalMux I__210 (
            .O(N__1458),
            .I(cntrZ0Z_0));
    LocalMux I__209 (
            .O(N__1455),
            .I(cntrZ0Z_0));
    CascadeMux I__208 (
            .O(N__1446),
            .I(BIT_47_i_o3_0_0_4_cascade_));
    CascadeMux I__207 (
            .O(N__1443),
            .I(N__1437));
    InMux I__206 (
            .O(N__1442),
            .I(N__1434));
    InMux I__205 (
            .O(N__1441),
            .I(N__1427));
    InMux I__204 (
            .O(N__1440),
            .I(N__1427));
    InMux I__203 (
            .O(N__1437),
            .I(N__1427));
    LocalMux I__202 (
            .O(N__1434),
            .I(N_27));
    LocalMux I__201 (
            .O(N__1427),
            .I(N_27));
    InMux I__200 (
            .O(N__1422),
            .I(N__1410));
    InMux I__199 (
            .O(N__1421),
            .I(N__1410));
    InMux I__198 (
            .O(N__1420),
            .I(N__1410));
    InMux I__197 (
            .O(N__1419),
            .I(N__1410));
    LocalMux I__196 (
            .O(N__1410),
            .I(N_45));
    InMux I__195 (
            .O(N__1407),
            .I(N__1402));
    InMux I__194 (
            .O(N__1406),
            .I(N__1399));
    InMux I__193 (
            .O(N__1405),
            .I(N__1396));
    LocalMux I__192 (
            .O(N__1402),
            .I(N_17));
    LocalMux I__191 (
            .O(N__1399),
            .I(N_17));
    LocalMux I__190 (
            .O(N__1396),
            .I(N_17));
    CascadeMux I__189 (
            .O(N__1389),
            .I(N_45_cascade_));
    CascadeMux I__188 (
            .O(N__1386),
            .I(N__1383));
    InMux I__187 (
            .O(N__1383),
            .I(N__1377));
    InMux I__186 (
            .O(N__1382),
            .I(N__1377));
    LocalMux I__185 (
            .O(N__1377),
            .I(N_30));
    InMux I__184 (
            .O(N__1374),
            .I(bfn_2_6_0_));
    InMux I__183 (
            .O(N__1371),
            .I(N__1364));
    InMux I__182 (
            .O(N__1370),
            .I(N__1361));
    InMux I__181 (
            .O(N__1369),
            .I(N__1356));
    InMux I__180 (
            .O(N__1368),
            .I(N__1356));
    InMux I__179 (
            .O(N__1367),
            .I(N__1353));
    LocalMux I__178 (
            .O(N__1364),
            .I(cntrZ0Z_1));
    LocalMux I__177 (
            .O(N__1361),
            .I(cntrZ0Z_1));
    LocalMux I__176 (
            .O(N__1356),
            .I(cntrZ0Z_1));
    LocalMux I__175 (
            .O(N__1353),
            .I(cntrZ0Z_1));
    InMux I__174 (
            .O(N__1344),
            .I(cntr_cry_0));
    InMux I__173 (
            .O(N__1341),
            .I(cntr_cry_1));
    InMux I__172 (
            .O(N__1338),
            .I(cntr_cry_2));
    InMux I__171 (
            .O(N__1335),
            .I(clk_div_2_cry_18));
    InMux I__170 (
            .O(N__1332),
            .I(N__1329));
    LocalMux I__169 (
            .O(N__1329),
            .I(BIT_47_0));
    IoInMux I__168 (
            .O(N__1326),
            .I(N__1323));
    LocalMux I__167 (
            .O(N__1323),
            .I(N__1320));
    Span4Mux_s2_v I__166 (
            .O(N__1320),
            .I(N__1317));
    Span4Mux_v I__165 (
            .O(N__1317),
            .I(N__1313));
    CascadeMux I__164 (
            .O(N__1316),
            .I(N__1310));
    Span4Mux_h I__163 (
            .O(N__1313),
            .I(N__1306));
    InMux I__162 (
            .O(N__1310),
            .I(N__1303));
    InMux I__161 (
            .O(N__1309),
            .I(N__1300));
    Odrv4 I__160 (
            .O(N__1306),
            .I(LED0_c));
    LocalMux I__159 (
            .O(N__1303),
            .I(LED0_c));
    LocalMux I__158 (
            .O(N__1300),
            .I(LED0_c));
    CascadeMux I__157 (
            .O(N__1293),
            .I(clk_div_RNIICCP5Z0Z_19_cascade_));
    InMux I__156 (
            .O(N__1290),
            .I(N__1287));
    LocalMux I__155 (
            .O(N__1287),
            .I(N_12_i));
    IoInMux I__154 (
            .O(N__1284),
            .I(N__1281));
    LocalMux I__153 (
            .O(N__1281),
            .I(N__1277));
    CascadeMux I__152 (
            .O(N__1280),
            .I(N__1274));
    Span4Mux_s2_v I__151 (
            .O(N__1277),
            .I(N__1270));
    InMux I__150 (
            .O(N__1274),
            .I(N__1267));
    InMux I__149 (
            .O(N__1273),
            .I(N__1264));
    Span4Mux_h I__148 (
            .O(N__1270),
            .I(N__1261));
    LocalMux I__147 (
            .O(N__1267),
            .I(N__1256));
    LocalMux I__146 (
            .O(N__1264),
            .I(N__1256));
    Odrv4 I__145 (
            .O(N__1261),
            .I(LED2_c));
    Odrv4 I__144 (
            .O(N__1256),
            .I(LED2_c));
    InMux I__143 (
            .O(N__1251),
            .I(N__1248));
    LocalMux I__142 (
            .O(N__1248),
            .I(N_14_i));
    IoInMux I__141 (
            .O(N__1245),
            .I(N__1242));
    LocalMux I__140 (
            .O(N__1242),
            .I(N__1238));
    CascadeMux I__139 (
            .O(N__1241),
            .I(N__1235));
    IoSpan4Mux I__138 (
            .O(N__1238),
            .I(N__1231));
    InMux I__137 (
            .O(N__1235),
            .I(N__1228));
    InMux I__136 (
            .O(N__1234),
            .I(N__1225));
    Odrv4 I__135 (
            .O(N__1231),
            .I(LED3_c));
    LocalMux I__134 (
            .O(N__1228),
            .I(LED3_c));
    LocalMux I__133 (
            .O(N__1225),
            .I(LED3_c));
    InMux I__132 (
            .O(N__1218),
            .I(N__1215));
    LocalMux I__131 (
            .O(N__1215),
            .I(N_6_i));
    IoInMux I__130 (
            .O(N__1212),
            .I(N__1209));
    LocalMux I__129 (
            .O(N__1209),
            .I(N__1206));
    Span4Mux_s2_v I__128 (
            .O(N__1206),
            .I(N__1202));
    CascadeMux I__127 (
            .O(N__1205),
            .I(N__1199));
    Span4Mux_v I__126 (
            .O(N__1202),
            .I(N__1195));
    InMux I__125 (
            .O(N__1199),
            .I(N__1192));
    InMux I__124 (
            .O(N__1198),
            .I(N__1189));
    Odrv4 I__123 (
            .O(N__1195),
            .I(LED4_c));
    LocalMux I__122 (
            .O(N__1192),
            .I(LED4_c));
    LocalMux I__121 (
            .O(N__1189),
            .I(LED4_c));
    InMux I__120 (
            .O(N__1182),
            .I(N__1179));
    LocalMux I__119 (
            .O(N__1179),
            .I(N_8_i));
    IoInMux I__118 (
            .O(N__1176),
            .I(N__1172));
    CascadeMux I__117 (
            .O(N__1175),
            .I(N__1169));
    LocalMux I__116 (
            .O(N__1172),
            .I(N__1165));
    InMux I__115 (
            .O(N__1169),
            .I(N__1162));
    InMux I__114 (
            .O(N__1168),
            .I(N__1159));
    Span4Mux_s0_h I__113 (
            .O(N__1165),
            .I(N__1152));
    LocalMux I__112 (
            .O(N__1162),
            .I(N__1152));
    LocalMux I__111 (
            .O(N__1159),
            .I(N__1152));
    Odrv4 I__110 (
            .O(N__1152),
            .I(LED5_c));
    CascadeMux I__109 (
            .O(N__1149),
            .I(N_17_cascade_));
    CascadeMux I__108 (
            .O(N__1146),
            .I(N_22_cascade_));
    CascadeMux I__107 (
            .O(N__1143),
            .I(N__1140));
    InMux I__106 (
            .O(N__1140),
            .I(N__1137));
    LocalMux I__105 (
            .O(N__1137),
            .I(BIT_47_0_a3_0_1_6));
    CascadeMux I__104 (
            .O(N__1134),
            .I(N__1131));
    InMux I__103 (
            .O(N__1131),
            .I(N__1125));
    InMux I__102 (
            .O(N__1130),
            .I(N__1125));
    LocalMux I__101 (
            .O(N__1125),
            .I(N__1122));
    Odrv4 I__100 (
            .O(N__1122),
            .I(N_31));
    CascadeMux I__99 (
            .O(N__1119),
            .I(BIT_47_0_a3_0_1_6_cascade_));
    defparam IN_MUX_bfv_1_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_8_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(clk_div_2_cry_8),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(clk_div_2_cry_16),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(clk_div_1_cry_8),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(clk_div_1_cry_16),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_2_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_6_0_));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam cntr_RNI1FK_0_LC_1_5_0.C_ON=1'b0;
    defparam cntr_RNI1FK_0_LC_1_5_0.SEQ_MODE=4'b0000;
    defparam cntr_RNI1FK_0_LC_1_5_0.LUT_INIT=16'b0001000100000000;
    LogicCell40 cntr_RNI1FK_0_LC_1_5_0 (
            .in0(N__1368),
            .in1(N__1470),
            .in2(_gnd_net_),
            .in3(N__2059),
            .lcout(BIT_47_0_a3_0_1_6),
            .ltout(BIT_47_0_a3_0_1_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNI9VF1_6_LC_1_5_1.C_ON=1'b0;
    defparam cntr_RNI9VF1_6_LC_1_5_1.SEQ_MODE=4'b0000;
    defparam cntr_RNI9VF1_6_LC_1_5_1.LUT_INIT=16'b0101000000100010;
    LogicCell40 cntr_RNI9VF1_6_LC_1_5_1 (
            .in0(N__1592),
            .in1(N__1405),
            .in2(N__1119),
            .in3(N__1510),
            .lcout(N_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNI3ND_2_LC_1_5_4.C_ON=1'b0;
    defparam cntr_RNI3ND_2_LC_1_5_4.SEQ_MODE=4'b0000;
    defparam cntr_RNI3ND_2_LC_1_5_4.LUT_INIT=16'b1111111100110011;
    LogicCell40 cntr_RNI3ND_2_LC_1_5_4 (
            .in0(_gnd_net_),
            .in1(N__2060),
            .in2(_gnd_net_),
            .in3(N__1543),
            .lcout(N_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNI8GR_0_LC_1_5_7.C_ON=1'b0;
    defparam cntr_RNI8GR_0_LC_1_5_7.SEQ_MODE=4'b0000;
    defparam cntr_RNI8GR_0_LC_1_5_7.LUT_INIT=16'b1101111111111111;
    LogicCell40 cntr_RNI8GR_0_LC_1_5_7 (
            .in0(N__1471),
            .in1(N__1509),
            .in2(N__1596),
            .in3(N__1369),
            .lcout(N_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNIVID_0_LC_1_6_0.C_ON=1'b0;
    defparam cntr_RNIVID_0_LC_1_6_0.SEQ_MODE=4'b0000;
    defparam cntr_RNIVID_0_LC_1_6_0.LUT_INIT=16'b0011001111111111;
    LogicCell40 cntr_RNIVID_0_LC_1_6_0 (
            .in0(_gnd_net_),
            .in1(N__1469),
            .in2(_gnd_net_),
            .in3(N__1367),
            .lcout(N_17),
            .ltout(N_17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNIC891_6_LC_1_6_1.C_ON=1'b0;
    defparam cntr_RNIC891_6_LC_1_6_1.SEQ_MODE=4'b0000;
    defparam cntr_RNIC891_6_LC_1_6_1.LUT_INIT=16'b1111110111111111;
    LogicCell40 cntr_RNIC891_6_LC_1_6_1 (
            .in0(N__1587),
            .in1(N__1505),
            .in2(N__1149),
            .in3(N__1419),
            .lcout(N_22),
            .ltout(N_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BIT_RNO_0_3_LC_1_6_2.C_ON=1'b0;
    defparam BIT_RNO_0_3_LC_1_6_2.SEQ_MODE=4'b0000;
    defparam BIT_RNO_0_3_LC_1_6_2.LUT_INIT=16'b1000000011000000;
    LogicCell40 BIT_RNO_0_3_LC_1_6_2 (
            .in0(N__1234),
            .in1(N__1442),
            .in2(N__1146),
            .in3(N__1382),
            .lcout(N_14_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNIE4G1_0_6_LC_1_6_3.C_ON=1'b0;
    defparam cntr_RNIE4G1_0_6_LC_1_6_3.SEQ_MODE=4'b0000;
    defparam cntr_RNIE4G1_0_6_LC_1_6_3.LUT_INIT=16'b0100000000000000;
    LogicCell40 cntr_RNIE4G1_0_6_LC_1_6_3 (
            .in0(N__1588),
            .in1(N__1506),
            .in2(N__1143),
            .in3(N__1420),
            .lcout(N_38),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BIT_RNO_0_0_LC_1_6_4.C_ON=1'b0;
    defparam BIT_RNO_0_0_LC_1_6_4.SEQ_MODE=4'b0000;
    defparam BIT_RNO_0_0_LC_1_6_4.LUT_INIT=16'b1010000010110011;
    LogicCell40 BIT_RNO_0_0_LC_1_6_4 (
            .in0(N__1309),
            .in1(N__1556),
            .in2(N__2028),
            .in3(N__1988),
            .lcout(BIT_47_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BIT_RNO_0_2_LC_1_6_5.C_ON=1'b0;
    defparam BIT_RNO_0_2_LC_1_6_5.SEQ_MODE=4'b0000;
    defparam BIT_RNO_0_2_LC_1_6_5.LUT_INIT=16'b0010101000111111;
    LogicCell40 BIT_RNO_0_2_LC_1_6_5 (
            .in0(N__1273),
            .in1(N__1421),
            .in2(N__1134),
            .in3(N__1440),
            .lcout(N_12_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BIT_RNO_0_5_LC_1_6_6.C_ON=1'b0;
    defparam BIT_RNO_0_5_LC_1_6_6.SEQ_MODE=4'b0000;
    defparam BIT_RNO_0_5_LC_1_6_6.LUT_INIT=16'b0111011100000111;
    LogicCell40 BIT_RNO_0_5_LC_1_6_6 (
            .in0(N__1422),
            .in1(N__1130),
            .in2(N__1443),
            .in3(N__1168),
            .lcout(N_8_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BIT_RNO_0_4_LC_1_6_7.C_ON=1'b0;
    defparam BIT_RNO_0_4_LC_1_6_7.SEQ_MODE=4'b0000;
    defparam BIT_RNO_0_4_LC_1_6_7.LUT_INIT=16'b1000101000000000;
    LogicCell40 BIT_RNO_0_4_LC_1_6_7 (
            .in0(N__2027),
            .in1(N__1198),
            .in2(N__1386),
            .in3(N__1441),
            .lcout(N_6_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BIT_0_LC_1_7_1.C_ON=1'b0;
    defparam BIT_0_LC_1_7_1.SEQ_MODE=4'b1000;
    defparam BIT_0_LC_1_7_1.LUT_INIT=16'b1111111011011100;
    LogicCell40 BIT_0_LC_1_7_1 (
            .in0(N__1804),
            .in1(N__1763),
            .in2(N__1316),
            .in3(N__1332),
            .lcout(LED0_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2262),
            .ce(),
            .sr(N__1709));
    defparam clk_div_RNIICCP5_19_LC_1_7_2.C_ON=1'b0;
    defparam clk_div_RNIICCP5_19_LC_1_7_2.SEQ_MODE=4'b0000;
    defparam clk_div_RNIICCP5_19_LC_1_7_2.LUT_INIT=16'b0011001100000000;
    LogicCell40 clk_div_RNIICCP5_19_LC_1_7_2 (
            .in0(_gnd_net_),
            .in1(N__2091),
            .in2(_gnd_net_),
            .in3(N__1879),
            .lcout(clk_div_RNIICCP5Z0Z_19),
            .ltout(clk_div_RNIICCP5Z0Z_19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BIT_1_LC_1_7_3.C_ON=1'b0;
    defparam BIT_1_LC_1_7_3.SEQ_MODE=4'b1000;
    defparam BIT_1_LC_1_7_3.LUT_INIT=16'b1111111110101100;
    LogicCell40 BIT_1_LC_1_7_3 (
            .in0(N__1938),
            .in1(N__1966),
            .in2(N__1293),
            .in3(N__1764),
            .lcout(LED1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2262),
            .ce(),
            .sr(N__1709));
    defparam BIT_2_LC_1_7_4.C_ON=1'b0;
    defparam BIT_2_LC_1_7_4.SEQ_MODE=4'b1000;
    defparam BIT_2_LC_1_7_4.LUT_INIT=16'b1111111010111010;
    LogicCell40 BIT_2_LC_1_7_4 (
            .in0(N__1761),
            .in1(N__1802),
            .in2(N__1280),
            .in3(N__1290),
            .lcout(LED2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2262),
            .ce(),
            .sr(N__1709));
    defparam BIT_3_LC_1_7_5.C_ON=1'b0;
    defparam BIT_3_LC_1_7_5.SEQ_MODE=4'b1000;
    defparam BIT_3_LC_1_7_5.LUT_INIT=16'b1111111011011100;
    LogicCell40 BIT_3_LC_1_7_5 (
            .in0(N__1805),
            .in1(N__1765),
            .in2(N__1241),
            .in3(N__1251),
            .lcout(LED3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2262),
            .ce(),
            .sr(N__1709));
    defparam BIT_4_LC_1_7_6.C_ON=1'b0;
    defparam BIT_4_LC_1_7_6.SEQ_MODE=4'b1000;
    defparam BIT_4_LC_1_7_6.LUT_INIT=16'b1111111010111010;
    LogicCell40 BIT_4_LC_1_7_6 (
            .in0(N__1762),
            .in1(N__1803),
            .in2(N__1205),
            .in3(N__1218),
            .lcout(LED4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2262),
            .ce(),
            .sr(N__1709));
    defparam BIT_5_LC_1_7_7.C_ON=1'b0;
    defparam BIT_5_LC_1_7_7.SEQ_MODE=4'b1000;
    defparam BIT_5_LC_1_7_7.LUT_INIT=16'b1111111011011100;
    LogicCell40 BIT_5_LC_1_7_7 (
            .in0(N__1806),
            .in1(N__1766),
            .in2(N__1175),
            .in3(N__1182),
            .lcout(LED5_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2262),
            .ce(),
            .sr(N__1709));
    defparam clk_div_RNI91U1_1_LC_1_8_0.C_ON=1'b1;
    defparam clk_div_RNI91U1_1_LC_1_8_0.SEQ_MODE=4'b0000;
    defparam clk_div_RNI91U1_1_LC_1_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNI91U1_1_LC_1_8_0 (
            .in0(_gnd_net_),
            .in1(N__1684),
            .in2(N__1664),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_8_0_),
            .carryout(clk_div_2_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIF3T2_2_LC_1_8_1.C_ON=1'b1;
    defparam clk_div_RNIF3T2_2_LC_1_8_1.SEQ_MODE=4'b0000;
    defparam clk_div_RNIF3T2_2_LC_1_8_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIF3T2_2_LC_1_8_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1638),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_1),
            .carryout(clk_div_2_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIM6S3_3_LC_1_8_2.C_ON=1'b1;
    defparam clk_div_RNIM6S3_3_LC_1_8_2.SEQ_MODE=4'b0000;
    defparam clk_div_RNIM6S3_3_LC_1_8_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIM6S3_3_LC_1_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__1620),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_2),
            .carryout(clk_div_2_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIUAR4_4_LC_1_8_3.C_ON=1'b1;
    defparam clk_div_RNIUAR4_4_LC_1_8_3.SEQ_MODE=4'b0000;
    defparam clk_div_RNIUAR4_4_LC_1_8_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIUAR4_4_LC_1_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2235),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_3),
            .carryout(clk_div_2_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNI7GQ5_5_LC_1_8_4.C_ON=1'b1;
    defparam clk_div_RNI7GQ5_5_LC_1_8_4.SEQ_MODE=4'b0000;
    defparam clk_div_RNI7GQ5_5_LC_1_8_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNI7GQ5_5_LC_1_8_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2217),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_4),
            .carryout(clk_div_2_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIHMP6_6_LC_1_8_5.C_ON=1'b1;
    defparam clk_div_RNIHMP6_6_LC_1_8_5.SEQ_MODE=4'b0000;
    defparam clk_div_RNIHMP6_6_LC_1_8_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIHMP6_6_LC_1_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2199),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_5),
            .carryout(clk_div_2_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNISTO7_7_LC_1_8_6.C_ON=1'b1;
    defparam clk_div_RNISTO7_7_LC_1_8_6.SEQ_MODE=4'b0000;
    defparam clk_div_RNISTO7_7_LC_1_8_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNISTO7_7_LC_1_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2181),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_6),
            .carryout(clk_div_2_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNI86O8_8_LC_1_8_7.C_ON=1'b1;
    defparam clk_div_RNI86O8_8_LC_1_8_7.SEQ_MODE=4'b0000;
    defparam clk_div_RNI86O8_8_LC_1_8_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNI86O8_8_LC_1_8_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2163),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_7),
            .carryout(clk_div_2_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNILFN9_9_LC_1_9_0.C_ON=1'b1;
    defparam clk_div_RNILFN9_9_LC_1_9_0.SEQ_MODE=4'b0000;
    defparam clk_div_RNILFN9_9_LC_1_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNILFN9_9_LC_1_9_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2145),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(clk_div_2_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIAAMP_10_LC_1_9_1.C_ON=1'b1;
    defparam clk_div_RNIAAMP_10_LC_1_9_1.SEQ_MODE=4'b0000;
    defparam clk_div_RNIAAMP_10_LC_1_9_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIAAMP_10_LC_1_9_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2127),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_9),
            .carryout(clk_div_2_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNI06L91_11_LC_1_9_2.C_ON=1'b1;
    defparam clk_div_RNI06L91_11_LC_1_9_2.SEQ_MODE=4'b0000;
    defparam clk_div_RNI06L91_11_LC_1_9_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNI06L91_11_LC_1_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2109),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_10),
            .carryout(clk_div_2_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIN2KP1_12_LC_1_9_3.C_ON=1'b1;
    defparam clk_div_RNIN2KP1_12_LC_1_9_3.SEQ_MODE=4'b0000;
    defparam clk_div_RNIN2KP1_12_LC_1_9_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIN2KP1_12_LC_1_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2391),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_11),
            .carryout(clk_div_2_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIF0J92_13_LC_1_9_4.C_ON=1'b1;
    defparam clk_div_RNIF0J92_13_LC_1_9_4.SEQ_MODE=4'b0000;
    defparam clk_div_RNIF0J92_13_LC_1_9_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIF0J92_13_LC_1_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2373),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_12),
            .carryout(clk_div_2_cry_13),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNI8VHP2_14_LC_1_9_5.C_ON=1'b1;
    defparam clk_div_RNI8VHP2_14_LC_1_9_5.SEQ_MODE=4'b0000;
    defparam clk_div_RNI8VHP2_14_LC_1_9_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNI8VHP2_14_LC_1_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2355),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_13),
            .carryout(clk_div_2_cry_14),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNI2VG93_15_LC_1_9_6.C_ON=1'b1;
    defparam clk_div_RNI2VG93_15_LC_1_9_6.SEQ_MODE=4'b0000;
    defparam clk_div_RNI2VG93_15_LC_1_9_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNI2VG93_15_LC_1_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2337),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_14),
            .carryout(clk_div_2_cry_15),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNITVFP3_16_LC_1_9_7.C_ON=1'b1;
    defparam clk_div_RNITVFP3_16_LC_1_9_7.SEQ_MODE=4'b0000;
    defparam clk_div_RNITVFP3_16_LC_1_9_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNITVFP3_16_LC_1_9_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2319),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_15),
            .carryout(clk_div_2_cry_16),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIP1F94_17_LC_1_10_0.C_ON=1'b1;
    defparam clk_div_RNIP1F94_17_LC_1_10_0.SEQ_MODE=4'b0000;
    defparam clk_div_RNIP1F94_17_LC_1_10_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIP1F94_17_LC_1_10_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2301),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(clk_div_2_cry_17),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIM4EP4_18_LC_1_10_1.C_ON=1'b1;
    defparam clk_div_RNIM4EP4_18_LC_1_10_1.SEQ_MODE=4'b0000;
    defparam clk_div_RNIM4EP4_18_LC_1_10_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIM4EP4_18_LC_1_10_1 (
            .in0(_gnd_net_),
            .in1(N__2279),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_17),
            .carryout(clk_div_2_cry_18),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIK8D95_19_LC_1_10_2.C_ON=1'b0;
    defparam clk_div_RNIK8D95_19_LC_1_10_2.SEQ_MODE=4'b0000;
    defparam clk_div_RNIK8D95_19_LC_1_10_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 clk_div_RNIK8D95_19_LC_1_10_2 (
            .in0(_gnd_net_),
            .in1(N__2075),
            .in2(_gnd_net_),
            .in3(N__1335),
            .lcout(clk_div_RNIK8D95Z0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_19_LC_1_10_7.C_ON=1'b0;
    defparam clk_div_19_LC_1_10_7.SEQ_MODE=4'b1000;
    defparam clk_div_19_LC_1_10_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 clk_div_19_LC_1_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1875),
            .lcout(clk_div_i_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2263),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNI6KK_2_LC_2_5_1.C_ON=1'b0;
    defparam cntr_RNI6KK_2_LC_2_5_1.SEQ_MODE=4'b0000;
    defparam cntr_RNI6KK_2_LC_2_5_1.LUT_INIT=16'b1111101011111111;
    LogicCell40 cntr_RNI6KK_2_LC_2_5_1 (
            .in0(N__1542),
            .in1(_gnd_net_),
            .in2(N__1931),
            .in3(N__2057),
            .lcout(),
            .ltout(BIT_47_i_o3_0_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNIE4G1_6_LC_2_5_2.C_ON=1'b0;
    defparam cntr_RNIE4G1_6_LC_2_5_2.SEQ_MODE=4'b0000;
    defparam cntr_RNIE4G1_6_LC_2_5_2.LUT_INIT=16'b1111111111111011;
    LogicCell40 cntr_RNIE4G1_6_LC_2_5_2 (
            .in0(N__1594),
            .in1(N__1507),
            .in2(N__1446),
            .in3(N__1407),
            .lcout(N_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNI4OD_2_LC_2_5_4.C_ON=1'b0;
    defparam cntr_RNI4OD_2_LC_2_5_4.SEQ_MODE=4'b0000;
    defparam cntr_RNI4OD_2_LC_2_5_4.LUT_INIT=16'b1100110000000000;
    LogicCell40 cntr_RNI4OD_2_LC_2_5_4 (
            .in0(_gnd_net_),
            .in1(N__1541),
            .in2(_gnd_net_),
            .in3(N__1922),
            .lcout(N_45),
            .ltout(N_45_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNI9591_3_LC_2_5_5.C_ON=1'b0;
    defparam cntr_RNI9591_3_LC_2_5_5.SEQ_MODE=4'b0000;
    defparam cntr_RNI9591_3_LC_2_5_5.LUT_INIT=16'b1111111111101111;
    LogicCell40 cntr_RNI9591_3_LC_2_5_5 (
            .in0(N__1508),
            .in1(N__1406),
            .in2(N__1389),
            .in3(N__2058),
            .lcout(N_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNI5PD_1_LC_2_5_7.C_ON=1'b0;
    defparam cntr_RNI5PD_1_LC_2_5_7.SEQ_MODE=4'b0000;
    defparam cntr_RNI5PD_1_LC_2_5_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 cntr_RNI5PD_1_LC_2_5_7 (
            .in0(_gnd_net_),
            .in1(N__1593),
            .in2(_gnd_net_),
            .in3(N__1370),
            .lcout(g0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_0_LC_2_6_0.C_ON=1'b1;
    defparam cntr_0_LC_2_6_0.SEQ_MODE=4'b1000;
    defparam cntr_0_LC_2_6_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_0_LC_2_6_0 (
            .in0(_gnd_net_),
            .in1(N__1473),
            .in2(_gnd_net_),
            .in3(N__1374),
            .lcout(cntrZ0Z_0),
            .ltout(),
            .carryin(bfn_2_6_0_),
            .carryout(cntr_cry_0),
            .clk(N__2267),
            .ce(N__1807),
            .sr(_gnd_net_));
    defparam cntr_1_LC_2_6_1.C_ON=1'b1;
    defparam cntr_1_LC_2_6_1.SEQ_MODE=4'b1000;
    defparam cntr_1_LC_2_6_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_1_LC_2_6_1 (
            .in0(_gnd_net_),
            .in1(N__1371),
            .in2(_gnd_net_),
            .in3(N__1344),
            .lcout(cntrZ0Z_1),
            .ltout(),
            .carryin(cntr_cry_0),
            .carryout(cntr_cry_1),
            .clk(N__2267),
            .ce(N__1807),
            .sr(_gnd_net_));
    defparam cntr_2_LC_2_6_2.C_ON=1'b1;
    defparam cntr_2_LC_2_6_2.SEQ_MODE=4'b1000;
    defparam cntr_2_LC_2_6_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_2_LC_2_6_2 (
            .in0(_gnd_net_),
            .in1(N__1545),
            .in2(_gnd_net_),
            .in3(N__1341),
            .lcout(cntrZ0Z_2),
            .ltout(),
            .carryin(cntr_cry_1),
            .carryout(cntr_cry_2),
            .clk(N__2267),
            .ce(N__1807),
            .sr(_gnd_net_));
    defparam cntr_3_LC_2_6_3.C_ON=1'b1;
    defparam cntr_3_LC_2_6_3.SEQ_MODE=4'b1000;
    defparam cntr_3_LC_2_6_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_3_LC_2_6_3 (
            .in0(_gnd_net_),
            .in1(N__2064),
            .in2(_gnd_net_),
            .in3(N__1338),
            .lcout(cntrZ0Z_3),
            .ltout(),
            .carryin(cntr_cry_2),
            .carryout(cntr_cry_3),
            .clk(N__2267),
            .ce(N__1807),
            .sr(_gnd_net_));
    defparam cntr_4_LC_2_6_4.C_ON=1'b1;
    defparam cntr_4_LC_2_6_4.SEQ_MODE=4'b1000;
    defparam cntr_4_LC_2_6_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_4_LC_2_6_4 (
            .in0(_gnd_net_),
            .in1(N__1930),
            .in2(_gnd_net_),
            .in3(N__1605),
            .lcout(cntrZ0Z_4),
            .ltout(),
            .carryin(cntr_cry_3),
            .carryout(cntr_cry_4),
            .clk(N__2267),
            .ce(N__1807),
            .sr(_gnd_net_));
    defparam cntr_5_LC_2_6_5.C_ON=1'b1;
    defparam cntr_5_LC_2_6_5.SEQ_MODE=4'b1000;
    defparam cntr_5_LC_2_6_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_5_LC_2_6_5 (
            .in0(_gnd_net_),
            .in1(N__1514),
            .in2(_gnd_net_),
            .in3(N__1602),
            .lcout(cntrZ0Z_5),
            .ltout(),
            .carryin(cntr_cry_4),
            .carryout(cntr_cry_5),
            .clk(N__2267),
            .ce(N__1807),
            .sr(_gnd_net_));
    defparam cntr_6_LC_2_6_6.C_ON=1'b0;
    defparam cntr_6_LC_2_6_6.SEQ_MODE=4'b1000;
    defparam cntr_6_LC_2_6_6.LUT_INIT=16'b0011001111001100;
    LogicCell40 cntr_6_LC_2_6_6 (
            .in0(_gnd_net_),
            .in1(N__1595),
            .in2(_gnd_net_),
            .in3(N__1599),
            .lcout(cntrZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2267),
            .ce(N__1807),
            .sr(_gnd_net_));
    defparam BIT_RNO_0_7_LC_2_7_0.C_ON=1'b0;
    defparam BIT_RNO_0_7_LC_2_7_0.SEQ_MODE=4'b0000;
    defparam BIT_RNO_0_7_LC_2_7_0.LUT_INIT=16'b1111000100010001;
    LogicCell40 BIT_RNO_0_7_LC_2_7_0 (
            .in0(N__1998),
            .in1(N__1560),
            .in2(N__1736),
            .in3(N__2023),
            .lcout(BIT_47_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_1_LC_2_7_1.C_ON=1'b0;
    defparam clk_div_1_LC_2_7_1.SEQ_MODE=4'b1000;
    defparam clk_div_1_LC_2_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 clk_div_1_LC_2_7_1 (
            .in0(_gnd_net_),
            .in1(N__1662),
            .in2(_gnd_net_),
            .in3(N__1688),
            .lcout(clk_divZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2264),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNI6KK_0_2_LC_2_7_2.C_ON=1'b0;
    defparam cntr_RNI6KK_0_2_LC_2_7_2.SEQ_MODE=4'b0000;
    defparam cntr_RNI6KK_0_2_LC_2_7_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 cntr_RNI6KK_0_2_LC_2_7_2 (
            .in0(N__1926),
            .in1(N__2061),
            .in2(_gnd_net_),
            .in3(N__1544),
            .lcout(N_21),
            .ltout(N_21_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BIT_RNO_0_6_LC_2_7_3.C_ON=1'b0;
    defparam BIT_RNO_0_6_LC_2_7_3.SEQ_MODE=4'b0000;
    defparam BIT_RNO_0_6_LC_2_7_3.LUT_INIT=16'b1111111110001010;
    LogicCell40 BIT_RNO_0_6_LC_2_7_3 (
            .in0(N__1832),
            .in1(N__1997),
            .in2(N__1518),
            .in3(N__1947),
            .lcout(BIT_47_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNI3NJG_19_LC_2_7_4.C_ON=1'b0;
    defparam clk_div_RNI3NJG_19_LC_2_7_4.SEQ_MODE=4'b0000;
    defparam clk_div_RNI3NJG_19_LC_2_7_4.LUT_INIT=16'b0000010000000000;
    LogicCell40 clk_div_RNI3NJG_19_LC_2_7_4 (
            .in0(N__2089),
            .in1(N__2062),
            .in2(N__1515),
            .in3(N__1472),
            .lcout(g0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_0_LC_2_7_5.C_ON=1'b0;
    defparam clk_div_0_LC_2_7_5.SEQ_MODE=4'b1000;
    defparam clk_div_0_LC_2_7_5.LUT_INIT=16'b0000000011111111;
    LogicCell40 clk_div_0_LC_2_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1663),
            .lcout(clk_divZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2264),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNI0HSQ5_19_LC_2_7_6.C_ON=1'b0;
    defparam clk_div_RNI0HSQ5_19_LC_2_7_6.SEQ_MODE=4'b0000;
    defparam clk_div_RNI0HSQ5_19_LC_2_7_6.LUT_INIT=16'b0000000001000000;
    LogicCell40 clk_div_RNI0HSQ5_19_LC_2_7_6 (
            .in0(N__2090),
            .in1(N__2063),
            .in2(N__1881),
            .in3(N__2022),
            .lcout(clk_div_RNI0HSQ5Z0Z_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BIT_RNO_0_1_LC_2_7_7.C_ON=1'b0;
    defparam BIT_RNO_0_1_LC_2_7_7.SEQ_MODE=4'b0000;
    defparam BIT_RNO_0_1_LC_2_7_7.LUT_INIT=16'b1111111111010000;
    LogicCell40 BIT_RNO_0_1_LC_2_7_7 (
            .in0(N__2004),
            .in1(N__1996),
            .in2(N__1976),
            .in3(N__1946),
            .lcout(BIT_47_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNIVLLQ5_4_LC_2_8_2.C_ON=1'b0;
    defparam cntr_RNIVLLQ5_4_LC_2_8_2.SEQ_MODE=4'b0000;
    defparam cntr_RNIVLLQ5_4_LC_2_8_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 cntr_RNIVLLQ5_4_LC_2_8_2 (
            .in0(N__1932),
            .in1(N__1899),
            .in2(N__1890),
            .in3(N__1880),
            .lcout(cntr_RNIVLLQ5Z0Z_4),
            .ltout(cntr_RNIVLLQ5Z0Z_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BIT_6_LC_2_8_3.C_ON=1'b0;
    defparam BIT_6_LC_2_8_3.SEQ_MODE=4'b1000;
    defparam BIT_6_LC_2_8_3.LUT_INIT=16'b1111111011110100;
    LogicCell40 BIT_6_LC_2_8_3 (
            .in0(N__1808),
            .in1(N__1828),
            .in2(N__1845),
            .in3(N__1842),
            .lcout(LED6_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2261),
            .ce(),
            .sr(N__1710));
    defparam BIT_7_LC_2_8_5.C_ON=1'b0;
    defparam BIT_7_LC_2_8_5.SEQ_MODE=4'b1000;
    defparam BIT_7_LC_2_8_5.LUT_INIT=16'b1111111111100100;
    LogicCell40 BIT_7_LC_2_8_5 (
            .in0(N__1809),
            .in1(N__1729),
            .in2(N__1776),
            .in3(N__1767),
            .lcout(LED7_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2261),
            .ce(),
            .sr(N__1710));
    defparam clk_div_1_cry_1_c_LC_2_9_0.C_ON=1'b1;
    defparam clk_div_1_cry_1_c_LC_2_9_0.SEQ_MODE=4'b0000;
    defparam clk_div_1_cry_1_c_LC_2_9_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_1_cry_1_c_LC_2_9_0 (
            .in0(_gnd_net_),
            .in1(N__1689),
            .in2(N__1668),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(clk_div_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_2_LC_2_9_1.C_ON=1'b1;
    defparam clk_div_2_LC_2_9_1.SEQ_MODE=4'b1000;
    defparam clk_div_2_LC_2_9_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_2_LC_2_9_1 (
            .in0(_gnd_net_),
            .in1(N__1637),
            .in2(_gnd_net_),
            .in3(N__1623),
            .lcout(clk_divZ0Z_2),
            .ltout(),
            .carryin(clk_div_1_cry_1),
            .carryout(clk_div_1_cry_2),
            .clk(N__2265),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_3_LC_2_9_2.C_ON=1'b1;
    defparam clk_div_3_LC_2_9_2.SEQ_MODE=4'b1000;
    defparam clk_div_3_LC_2_9_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_3_LC_2_9_2 (
            .in0(_gnd_net_),
            .in1(N__1619),
            .in2(_gnd_net_),
            .in3(N__2238),
            .lcout(clk_divZ0Z_3),
            .ltout(),
            .carryin(clk_div_1_cry_2),
            .carryout(clk_div_1_cry_3),
            .clk(N__2265),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_4_LC_2_9_3.C_ON=1'b1;
    defparam clk_div_4_LC_2_9_3.SEQ_MODE=4'b1000;
    defparam clk_div_4_LC_2_9_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_4_LC_2_9_3 (
            .in0(_gnd_net_),
            .in1(N__2234),
            .in2(_gnd_net_),
            .in3(N__2220),
            .lcout(clk_divZ0Z_4),
            .ltout(),
            .carryin(clk_div_1_cry_3),
            .carryout(clk_div_1_cry_4),
            .clk(N__2265),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_5_LC_2_9_4.C_ON=1'b1;
    defparam clk_div_5_LC_2_9_4.SEQ_MODE=4'b1000;
    defparam clk_div_5_LC_2_9_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_5_LC_2_9_4 (
            .in0(_gnd_net_),
            .in1(N__2216),
            .in2(_gnd_net_),
            .in3(N__2202),
            .lcout(clk_divZ0Z_5),
            .ltout(),
            .carryin(clk_div_1_cry_4),
            .carryout(clk_div_1_cry_5),
            .clk(N__2265),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_6_LC_2_9_5.C_ON=1'b1;
    defparam clk_div_6_LC_2_9_5.SEQ_MODE=4'b1000;
    defparam clk_div_6_LC_2_9_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_6_LC_2_9_5 (
            .in0(_gnd_net_),
            .in1(N__2198),
            .in2(_gnd_net_),
            .in3(N__2184),
            .lcout(clk_divZ0Z_6),
            .ltout(),
            .carryin(clk_div_1_cry_5),
            .carryout(clk_div_1_cry_6),
            .clk(N__2265),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_7_LC_2_9_6.C_ON=1'b1;
    defparam clk_div_7_LC_2_9_6.SEQ_MODE=4'b1000;
    defparam clk_div_7_LC_2_9_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_7_LC_2_9_6 (
            .in0(_gnd_net_),
            .in1(N__2180),
            .in2(_gnd_net_),
            .in3(N__2166),
            .lcout(clk_divZ0Z_7),
            .ltout(),
            .carryin(clk_div_1_cry_6),
            .carryout(clk_div_1_cry_7),
            .clk(N__2265),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_8_LC_2_9_7.C_ON=1'b1;
    defparam clk_div_8_LC_2_9_7.SEQ_MODE=4'b1000;
    defparam clk_div_8_LC_2_9_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_8_LC_2_9_7 (
            .in0(_gnd_net_),
            .in1(N__2162),
            .in2(_gnd_net_),
            .in3(N__2148),
            .lcout(clk_divZ0Z_8),
            .ltout(),
            .carryin(clk_div_1_cry_7),
            .carryout(clk_div_1_cry_8),
            .clk(N__2265),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_9_LC_2_10_0.C_ON=1'b1;
    defparam clk_div_9_LC_2_10_0.SEQ_MODE=4'b1000;
    defparam clk_div_9_LC_2_10_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_9_LC_2_10_0 (
            .in0(_gnd_net_),
            .in1(N__2144),
            .in2(_gnd_net_),
            .in3(N__2130),
            .lcout(clk_divZ0Z_9),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(clk_div_1_cry_9),
            .clk(N__2266),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_10_LC_2_10_1.C_ON=1'b1;
    defparam clk_div_10_LC_2_10_1.SEQ_MODE=4'b1000;
    defparam clk_div_10_LC_2_10_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_10_LC_2_10_1 (
            .in0(_gnd_net_),
            .in1(N__2126),
            .in2(_gnd_net_),
            .in3(N__2112),
            .lcout(clk_divZ0Z_10),
            .ltout(),
            .carryin(clk_div_1_cry_9),
            .carryout(clk_div_1_cry_10),
            .clk(N__2266),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_11_LC_2_10_2.C_ON=1'b1;
    defparam clk_div_11_LC_2_10_2.SEQ_MODE=4'b1000;
    defparam clk_div_11_LC_2_10_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_11_LC_2_10_2 (
            .in0(_gnd_net_),
            .in1(N__2108),
            .in2(_gnd_net_),
            .in3(N__2094),
            .lcout(clk_divZ0Z_11),
            .ltout(),
            .carryin(clk_div_1_cry_10),
            .carryout(clk_div_1_cry_11),
            .clk(N__2266),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_12_LC_2_10_3.C_ON=1'b1;
    defparam clk_div_12_LC_2_10_3.SEQ_MODE=4'b1000;
    defparam clk_div_12_LC_2_10_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_12_LC_2_10_3 (
            .in0(_gnd_net_),
            .in1(N__2390),
            .in2(_gnd_net_),
            .in3(N__2376),
            .lcout(clk_divZ0Z_12),
            .ltout(),
            .carryin(clk_div_1_cry_11),
            .carryout(clk_div_1_cry_12),
            .clk(N__2266),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_13_LC_2_10_4.C_ON=1'b1;
    defparam clk_div_13_LC_2_10_4.SEQ_MODE=4'b1000;
    defparam clk_div_13_LC_2_10_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_13_LC_2_10_4 (
            .in0(_gnd_net_),
            .in1(N__2372),
            .in2(_gnd_net_),
            .in3(N__2358),
            .lcout(clk_divZ0Z_13),
            .ltout(),
            .carryin(clk_div_1_cry_12),
            .carryout(clk_div_1_cry_13),
            .clk(N__2266),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_14_LC_2_10_5.C_ON=1'b1;
    defparam clk_div_14_LC_2_10_5.SEQ_MODE=4'b1000;
    defparam clk_div_14_LC_2_10_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_14_LC_2_10_5 (
            .in0(_gnd_net_),
            .in1(N__2354),
            .in2(_gnd_net_),
            .in3(N__2340),
            .lcout(clk_divZ0Z_14),
            .ltout(),
            .carryin(clk_div_1_cry_13),
            .carryout(clk_div_1_cry_14),
            .clk(N__2266),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_15_LC_2_10_6.C_ON=1'b1;
    defparam clk_div_15_LC_2_10_6.SEQ_MODE=4'b1000;
    defparam clk_div_15_LC_2_10_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_15_LC_2_10_6 (
            .in0(_gnd_net_),
            .in1(N__2336),
            .in2(_gnd_net_),
            .in3(N__2322),
            .lcout(clk_divZ0Z_15),
            .ltout(),
            .carryin(clk_div_1_cry_14),
            .carryout(clk_div_1_cry_15),
            .clk(N__2266),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_16_LC_2_10_7.C_ON=1'b1;
    defparam clk_div_16_LC_2_10_7.SEQ_MODE=4'b1000;
    defparam clk_div_16_LC_2_10_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_16_LC_2_10_7 (
            .in0(_gnd_net_),
            .in1(N__2318),
            .in2(_gnd_net_),
            .in3(N__2304),
            .lcout(clk_divZ0Z_16),
            .ltout(),
            .carryin(clk_div_1_cry_15),
            .carryout(clk_div_1_cry_16),
            .clk(N__2266),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_17_LC_2_11_0.C_ON=1'b1;
    defparam clk_div_17_LC_2_11_0.SEQ_MODE=4'b1000;
    defparam clk_div_17_LC_2_11_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_17_LC_2_11_0 (
            .in0(_gnd_net_),
            .in1(N__2300),
            .in2(_gnd_net_),
            .in3(N__2286),
            .lcout(clk_divZ0Z_17),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(clk_div_1_cry_17),
            .clk(N__2268),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_18_LC_2_11_1.C_ON=1'b0;
    defparam clk_div_18_LC_2_11_1.SEQ_MODE=4'b1000;
    defparam clk_div_18_LC_2_11_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 clk_div_18_LC_2_11_1 (
            .in0(_gnd_net_),
            .in1(N__2280),
            .in2(_gnd_net_),
            .in3(N__2283),
            .lcout(clk_divZ0Z_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2268),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
