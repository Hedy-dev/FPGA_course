-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jul 13 2021 15:22:48

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    LED5 : out std_logic;
    LED1 : out std_logic;
    LED6 : out std_logic;
    LED4 : out std_logic;
    LED2 : out std_logic;
    LED0 : out std_logic;
    CLK : in std_logic;
    LED7 : out std_logic;
    LED3 : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__2484\ : std_logic;
signal \N__2483\ : std_logic;
signal \N__2482\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2471\ : std_logic;
signal \N__2464\ : std_logic;
signal \N__2463\ : std_logic;
signal \N__2462\ : std_logic;
signal \N__2455\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2445\ : std_logic;
signal \N__2444\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2436\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2426\ : std_logic;
signal \N__2419\ : std_logic;
signal \N__2418\ : std_logic;
signal \N__2417\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2408\ : std_logic;
signal \N__2391\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2384\ : std_logic;
signal \N__2381\ : std_logic;
signal \N__2376\ : std_logic;
signal \N__2373\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2369\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2358\ : std_logic;
signal \N__2355\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2340\ : std_logic;
signal \N__2337\ : std_logic;
signal \N__2336\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2322\ : std_logic;
signal \N__2319\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2304\ : std_logic;
signal \N__2301\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2294\ : std_logic;
signal \N__2291\ : std_logic;
signal \N__2286\ : std_logic;
signal \N__2283\ : std_logic;
signal \N__2280\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2268\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2266\ : std_logic;
signal \N__2265\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2263\ : std_logic;
signal \N__2262\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2244\ : std_logic;
signal \N__2241\ : std_logic;
signal \N__2238\ : std_logic;
signal \N__2235\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2228\ : std_logic;
signal \N__2225\ : std_logic;
signal \N__2220\ : std_logic;
signal \N__2217\ : std_logic;
signal \N__2216\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2207\ : std_logic;
signal \N__2202\ : std_logic;
signal \N__2199\ : std_logic;
signal \N__2198\ : std_logic;
signal \N__2195\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2184\ : std_logic;
signal \N__2181\ : std_logic;
signal \N__2180\ : std_logic;
signal \N__2177\ : std_logic;
signal \N__2174\ : std_logic;
signal \N__2171\ : std_logic;
signal \N__2166\ : std_logic;
signal \N__2163\ : std_logic;
signal \N__2162\ : std_logic;
signal \N__2159\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2153\ : std_logic;
signal \N__2148\ : std_logic;
signal \N__2145\ : std_logic;
signal \N__2144\ : std_logic;
signal \N__2141\ : std_logic;
signal \N__2138\ : std_logic;
signal \N__2135\ : std_logic;
signal \N__2130\ : std_logic;
signal \N__2127\ : std_logic;
signal \N__2126\ : std_logic;
signal \N__2123\ : std_logic;
signal \N__2120\ : std_logic;
signal \N__2117\ : std_logic;
signal \N__2112\ : std_logic;
signal \N__2109\ : std_logic;
signal \N__2108\ : std_logic;
signal \N__2105\ : std_logic;
signal \N__2102\ : std_logic;
signal \N__2099\ : std_logic;
signal \N__2094\ : std_logic;
signal \N__2091\ : std_logic;
signal \N__2090\ : std_logic;
signal \N__2089\ : std_logic;
signal \N__2086\ : std_logic;
signal \N__2081\ : std_logic;
signal \N__2076\ : std_logic;
signal \N__2075\ : std_logic;
signal \N__2072\ : std_logic;
signal \N__2069\ : std_logic;
signal \N__2064\ : std_logic;
signal \N__2063\ : std_logic;
signal \N__2062\ : std_logic;
signal \N__2061\ : std_logic;
signal \N__2060\ : std_logic;
signal \N__2059\ : std_logic;
signal \N__2058\ : std_logic;
signal \N__2057\ : std_logic;
signal \N__2054\ : std_logic;
signal \N__2047\ : std_logic;
signal \N__2042\ : std_logic;
signal \N__2037\ : std_logic;
signal \N__2028\ : std_logic;
signal \N__2027\ : std_logic;
signal \N__2024\ : std_logic;
signal \N__2023\ : std_logic;
signal \N__2022\ : std_logic;
signal \N__2019\ : std_logic;
signal \N__2016\ : std_logic;
signal \N__2011\ : std_logic;
signal \N__2004\ : std_logic;
signal \N__2001\ : std_logic;
signal \N__1998\ : std_logic;
signal \N__1997\ : std_logic;
signal \N__1996\ : std_logic;
signal \N__1989\ : std_logic;
signal \N__1988\ : std_logic;
signal \N__1985\ : std_logic;
signal \N__1982\ : std_logic;
signal \N__1977\ : std_logic;
signal \N__1976\ : std_logic;
signal \N__1973\ : std_logic;
signal \N__1970\ : std_logic;
signal \N__1967\ : std_logic;
signal \N__1966\ : std_logic;
signal \N__1963\ : std_logic;
signal \N__1960\ : std_logic;
signal \N__1957\ : std_logic;
signal \N__1954\ : std_logic;
signal \N__1947\ : std_logic;
signal \N__1946\ : std_logic;
signal \N__1941\ : std_logic;
signal \N__1938\ : std_logic;
signal \N__1935\ : std_logic;
signal \N__1932\ : std_logic;
signal \N__1931\ : std_logic;
signal \N__1930\ : std_logic;
signal \N__1927\ : std_logic;
signal \N__1926\ : std_logic;
signal \N__1923\ : std_logic;
signal \N__1922\ : std_logic;
signal \N__1919\ : std_logic;
signal \N__1916\ : std_logic;
signal \N__1913\ : std_logic;
signal \N__1908\ : std_logic;
signal \N__1899\ : std_logic;
signal \N__1896\ : std_logic;
signal \N__1893\ : std_logic;
signal \N__1890\ : std_logic;
signal \N__1887\ : std_logic;
signal \N__1884\ : std_logic;
signal \N__1881\ : std_logic;
signal \N__1880\ : std_logic;
signal \N__1879\ : std_logic;
signal \N__1876\ : std_logic;
signal \N__1875\ : std_logic;
signal \N__1872\ : std_logic;
signal \N__1869\ : std_logic;
signal \N__1866\ : std_logic;
signal \N__1863\ : std_logic;
signal \N__1860\ : std_logic;
signal \N__1857\ : std_logic;
signal \N__1854\ : std_logic;
signal \N__1845\ : std_logic;
signal \N__1842\ : std_logic;
signal \N__1839\ : std_logic;
signal \N__1836\ : std_logic;
signal \N__1833\ : std_logic;
signal \N__1832\ : std_logic;
signal \N__1829\ : std_logic;
signal \N__1828\ : std_logic;
signal \N__1825\ : std_logic;
signal \N__1822\ : std_logic;
signal \N__1819\ : std_logic;
signal \N__1816\ : std_logic;
signal \N__1809\ : std_logic;
signal \N__1808\ : std_logic;
signal \N__1807\ : std_logic;
signal \N__1806\ : std_logic;
signal \N__1805\ : std_logic;
signal \N__1804\ : std_logic;
signal \N__1803\ : std_logic;
signal \N__1802\ : std_logic;
signal \N__1797\ : std_logic;
signal \N__1794\ : std_logic;
signal \N__1783\ : std_logic;
signal \N__1776\ : std_logic;
signal \N__1773\ : std_logic;
signal \N__1770\ : std_logic;
signal \N__1767\ : std_logic;
signal \N__1766\ : std_logic;
signal \N__1765\ : std_logic;
signal \N__1764\ : std_logic;
signal \N__1763\ : std_logic;
signal \N__1762\ : std_logic;
signal \N__1761\ : std_logic;
signal \N__1758\ : std_logic;
signal \N__1745\ : std_logic;
signal \N__1740\ : std_logic;
signal \N__1737\ : std_logic;
signal \N__1736\ : std_logic;
signal \N__1733\ : std_logic;
signal \N__1730\ : std_logic;
signal \N__1729\ : std_logic;
signal \N__1726\ : std_logic;
signal \N__1723\ : std_logic;
signal \N__1720\ : std_logic;
signal \N__1715\ : std_logic;
signal \N__1710\ : std_logic;
signal \N__1709\ : std_logic;
signal \N__1706\ : std_logic;
signal \N__1703\ : std_logic;
signal \N__1700\ : std_logic;
signal \N__1697\ : std_logic;
signal \N__1694\ : std_logic;
signal \N__1689\ : std_logic;
signal \N__1688\ : std_logic;
signal \N__1685\ : std_logic;
signal \N__1684\ : std_logic;
signal \N__1681\ : std_logic;
signal \N__1678\ : std_logic;
signal \N__1675\ : std_logic;
signal \N__1668\ : std_logic;
signal \N__1665\ : std_logic;
signal \N__1664\ : std_logic;
signal \N__1663\ : std_logic;
signal \N__1662\ : std_logic;
signal \N__1659\ : std_logic;
signal \N__1656\ : std_logic;
signal \N__1651\ : std_logic;
signal \N__1648\ : std_logic;
signal \N__1645\ : std_logic;
signal \N__1638\ : std_logic;
signal \N__1637\ : std_logic;
signal \N__1634\ : std_logic;
signal \N__1631\ : std_logic;
signal \N__1628\ : std_logic;
signal \N__1623\ : std_logic;
signal \N__1620\ : std_logic;
signal \N__1619\ : std_logic;
signal \N__1616\ : std_logic;
signal \N__1613\ : std_logic;
signal \N__1610\ : std_logic;
signal \N__1605\ : std_logic;
signal \N__1602\ : std_logic;
signal \N__1599\ : std_logic;
signal \N__1596\ : std_logic;
signal \N__1595\ : std_logic;
signal \N__1594\ : std_logic;
signal \N__1593\ : std_logic;
signal \N__1592\ : std_logic;
signal \N__1589\ : std_logic;
signal \N__1588\ : std_logic;
signal \N__1587\ : std_logic;
signal \N__1584\ : std_logic;
signal \N__1579\ : std_logic;
signal \N__1574\ : std_logic;
signal \N__1569\ : std_logic;
signal \N__1560\ : std_logic;
signal \N__1557\ : std_logic;
signal \N__1556\ : std_logic;
signal \N__1553\ : std_logic;
signal \N__1550\ : std_logic;
signal \N__1545\ : std_logic;
signal \N__1544\ : std_logic;
signal \N__1543\ : std_logic;
signal \N__1542\ : std_logic;
signal \N__1541\ : std_logic;
signal \N__1538\ : std_logic;
signal \N__1535\ : std_logic;
signal \N__1532\ : std_logic;
signal \N__1527\ : std_logic;
signal \N__1518\ : std_logic;
signal \N__1515\ : std_logic;
signal \N__1514\ : std_logic;
signal \N__1511\ : std_logic;
signal \N__1510\ : std_logic;
signal \N__1509\ : std_logic;
signal \N__1508\ : std_logic;
signal \N__1507\ : std_logic;
signal \N__1506\ : std_logic;
signal \N__1505\ : std_logic;
signal \N__1502\ : std_logic;
signal \N__1499\ : std_logic;
signal \N__1494\ : std_logic;
signal \N__1489\ : std_logic;
signal \N__1484\ : std_logic;
signal \N__1473\ : std_logic;
signal \N__1472\ : std_logic;
signal \N__1471\ : std_logic;
signal \N__1470\ : std_logic;
signal \N__1469\ : std_logic;
signal \N__1466\ : std_logic;
signal \N__1463\ : std_logic;
signal \N__1458\ : std_logic;
signal \N__1455\ : std_logic;
signal \N__1446\ : std_logic;
signal \N__1443\ : std_logic;
signal \N__1442\ : std_logic;
signal \N__1441\ : std_logic;
signal \N__1440\ : std_logic;
signal \N__1437\ : std_logic;
signal \N__1434\ : std_logic;
signal \N__1427\ : std_logic;
signal \N__1422\ : std_logic;
signal \N__1421\ : std_logic;
signal \N__1420\ : std_logic;
signal \N__1419\ : std_logic;
signal \N__1410\ : std_logic;
signal \N__1407\ : std_logic;
signal \N__1406\ : std_logic;
signal \N__1405\ : std_logic;
signal \N__1402\ : std_logic;
signal \N__1399\ : std_logic;
signal \N__1396\ : std_logic;
signal \N__1389\ : std_logic;
signal \N__1386\ : std_logic;
signal \N__1383\ : std_logic;
signal \N__1382\ : std_logic;
signal \N__1377\ : std_logic;
signal \N__1374\ : std_logic;
signal \N__1371\ : std_logic;
signal \N__1370\ : std_logic;
signal \N__1369\ : std_logic;
signal \N__1368\ : std_logic;
signal \N__1367\ : std_logic;
signal \N__1364\ : std_logic;
signal \N__1361\ : std_logic;
signal \N__1356\ : std_logic;
signal \N__1353\ : std_logic;
signal \N__1344\ : std_logic;
signal \N__1341\ : std_logic;
signal \N__1338\ : std_logic;
signal \N__1335\ : std_logic;
signal \N__1332\ : std_logic;
signal \N__1329\ : std_logic;
signal \N__1326\ : std_logic;
signal \N__1323\ : std_logic;
signal \N__1320\ : std_logic;
signal \N__1317\ : std_logic;
signal \N__1316\ : std_logic;
signal \N__1313\ : std_logic;
signal \N__1310\ : std_logic;
signal \N__1309\ : std_logic;
signal \N__1306\ : std_logic;
signal \N__1303\ : std_logic;
signal \N__1300\ : std_logic;
signal \N__1293\ : std_logic;
signal \N__1290\ : std_logic;
signal \N__1287\ : std_logic;
signal \N__1284\ : std_logic;
signal \N__1281\ : std_logic;
signal \N__1280\ : std_logic;
signal \N__1277\ : std_logic;
signal \N__1274\ : std_logic;
signal \N__1273\ : std_logic;
signal \N__1270\ : std_logic;
signal \N__1267\ : std_logic;
signal \N__1264\ : std_logic;
signal \N__1261\ : std_logic;
signal \N__1256\ : std_logic;
signal \N__1251\ : std_logic;
signal \N__1248\ : std_logic;
signal \N__1245\ : std_logic;
signal \N__1242\ : std_logic;
signal \N__1241\ : std_logic;
signal \N__1238\ : std_logic;
signal \N__1235\ : std_logic;
signal \N__1234\ : std_logic;
signal \N__1231\ : std_logic;
signal \N__1228\ : std_logic;
signal \N__1225\ : std_logic;
signal \N__1218\ : std_logic;
signal \N__1215\ : std_logic;
signal \N__1212\ : std_logic;
signal \N__1209\ : std_logic;
signal \N__1206\ : std_logic;
signal \N__1205\ : std_logic;
signal \N__1202\ : std_logic;
signal \N__1199\ : std_logic;
signal \N__1198\ : std_logic;
signal \N__1195\ : std_logic;
signal \N__1192\ : std_logic;
signal \N__1189\ : std_logic;
signal \N__1182\ : std_logic;
signal \N__1179\ : std_logic;
signal \N__1176\ : std_logic;
signal \N__1175\ : std_logic;
signal \N__1172\ : std_logic;
signal \N__1169\ : std_logic;
signal \N__1168\ : std_logic;
signal \N__1165\ : std_logic;
signal \N__1162\ : std_logic;
signal \N__1159\ : std_logic;
signal \N__1152\ : std_logic;
signal \N__1149\ : std_logic;
signal \N__1146\ : std_logic;
signal \N__1143\ : std_logic;
signal \N__1140\ : std_logic;
signal \N__1137\ : std_logic;
signal \N__1134\ : std_logic;
signal \N__1131\ : std_logic;
signal \N__1130\ : std_logic;
signal \N__1125\ : std_logic;
signal \N__1122\ : std_logic;
signal \N__1119\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \BIT_47_0_a3_0_1_6_cascade_\ : std_logic;
signal \N_17_cascade_\ : std_logic;
signal \N_22_cascade_\ : std_logic;
signal \BIT_47_0_a3_0_1_6\ : std_logic;
signal \N_31\ : std_logic;
signal \BIT_47_0\ : std_logic;
signal \LED0_c\ : std_logic;
signal \clk_div_RNIICCP5Z0Z_19_cascade_\ : std_logic;
signal \N_12_i\ : std_logic;
signal \LED2_c\ : std_logic;
signal \N_14_i\ : std_logic;
signal \LED3_c\ : std_logic;
signal \N_6_i\ : std_logic;
signal \LED4_c\ : std_logic;
signal \N_8_i\ : std_logic;
signal \LED5_c\ : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal clk_div_2_cry_1 : std_logic;
signal clk_div_2_cry_2 : std_logic;
signal clk_div_2_cry_3 : std_logic;
signal clk_div_2_cry_4 : std_logic;
signal clk_div_2_cry_5 : std_logic;
signal clk_div_2_cry_6 : std_logic;
signal clk_div_2_cry_7 : std_logic;
signal clk_div_2_cry_8 : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal clk_div_2_cry_9 : std_logic;
signal clk_div_2_cry_10 : std_logic;
signal clk_div_2_cry_11 : std_logic;
signal clk_div_2_cry_12 : std_logic;
signal clk_div_2_cry_13 : std_logic;
signal clk_div_2_cry_14 : std_logic;
signal clk_div_2_cry_15 : std_logic;
signal clk_div_2_cry_16 : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal clk_div_2_cry_17 : std_logic;
signal clk_div_2_cry_18 : std_logic;
signal \BIT_47_i_o3_0_0_4_cascade_\ : std_logic;
signal \N_27\ : std_logic;
signal \N_45\ : std_logic;
signal \N_17\ : std_logic;
signal \N_45_cascade_\ : std_logic;
signal \N_30\ : std_logic;
signal \bfn_2_6_0_\ : std_logic;
signal \cntrZ0Z_1\ : std_logic;
signal cntr_cry_0 : std_logic;
signal cntr_cry_1 : std_logic;
signal cntr_cry_2 : std_logic;
signal cntr_cry_3 : std_logic;
signal cntr_cry_4 : std_logic;
signal cntr_cry_5 : std_logic;
signal \cntrZ0Z_6\ : std_logic;
signal \N_23\ : std_logic;
signal \cntrZ0Z_2\ : std_logic;
signal \N_21_cascade_\ : std_logic;
signal \cntrZ0Z_5\ : std_logic;
signal \cntrZ0Z_0\ : std_logic;
signal clk_div_i_19 : std_logic;
signal \cntrZ0Z_3\ : std_logic;
signal \N_22\ : std_logic;
signal \N_21\ : std_logic;
signal \N_19\ : std_logic;
signal \LED1_c\ : std_logic;
signal \N_38\ : std_logic;
signal \BIT_47_1\ : std_logic;
signal \cntrZ0Z_4\ : std_logic;
signal g0_0 : std_logic;
signal g0_4 : std_logic;
signal \clk_div_RNIK8D95Z0Z_19\ : std_logic;
signal \cntr_RNIVLLQ5Z0Z_4_cascade_\ : std_logic;
signal \BIT_47_6\ : std_logic;
signal \LED6_c\ : std_logic;
signal \clk_div_RNIICCP5Z0Z_19\ : std_logic;
signal \BIT_47_7\ : std_logic;
signal \cntr_RNIVLLQ5Z0Z_4\ : std_logic;
signal \LED7_c\ : std_logic;
signal \clk_div_RNI0HSQ5Z0Z_19\ : std_logic;
signal \clk_divZ0Z_1\ : std_logic;
signal \clk_divZ0Z_0\ : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal \clk_divZ0Z_2\ : std_logic;
signal clk_div_1_cry_1 : std_logic;
signal \clk_divZ0Z_3\ : std_logic;
signal clk_div_1_cry_2 : std_logic;
signal \clk_divZ0Z_4\ : std_logic;
signal clk_div_1_cry_3 : std_logic;
signal \clk_divZ0Z_5\ : std_logic;
signal clk_div_1_cry_4 : std_logic;
signal \clk_divZ0Z_6\ : std_logic;
signal clk_div_1_cry_5 : std_logic;
signal \clk_divZ0Z_7\ : std_logic;
signal clk_div_1_cry_6 : std_logic;
signal \clk_divZ0Z_8\ : std_logic;
signal clk_div_1_cry_7 : std_logic;
signal clk_div_1_cry_8 : std_logic;
signal \clk_divZ0Z_9\ : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal \clk_divZ0Z_10\ : std_logic;
signal clk_div_1_cry_9 : std_logic;
signal \clk_divZ0Z_11\ : std_logic;
signal clk_div_1_cry_10 : std_logic;
signal \clk_divZ0Z_12\ : std_logic;
signal clk_div_1_cry_11 : std_logic;
signal \clk_divZ0Z_13\ : std_logic;
signal clk_div_1_cry_12 : std_logic;
signal \clk_divZ0Z_14\ : std_logic;
signal clk_div_1_cry_13 : std_logic;
signal \clk_divZ0Z_15\ : std_logic;
signal clk_div_1_cry_14 : std_logic;
signal \clk_divZ0Z_16\ : std_logic;
signal clk_div_1_cry_15 : std_logic;
signal clk_div_1_cry_16 : std_logic;
signal \clk_divZ0Z_17\ : std_logic;
signal \bfn_2_11_0_\ : std_logic;
signal clk_div_1_cry_17 : std_logic;
signal \clk_divZ0Z_18\ : std_logic;
signal \CLK_0_c_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK_wire\ : std_logic;
signal \LED4_wire\ : std_logic;
signal \LED2_wire\ : std_logic;
signal \LED0_wire\ : std_logic;
signal \LED6_wire\ : std_logic;
signal \LED3_wire\ : std_logic;
signal \LED7_wire\ : std_logic;
signal \LED1_wire\ : std_logic;
signal \LED5_wire\ : std_logic;

begin
    \CLK_wire\ <= CLK;
    LED4 <= \LED4_wire\;
    LED2 <= \LED2_wire\;
    LED0 <= \LED0_wire\;
    LED6 <= \LED6_wire\;
    LED3 <= \LED3_wire\;
    LED7 <= \LED7_wire\;
    LED1 <= \LED1_wire\;
    LED5 <= \LED5_wire\;

    \CLK_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__2482\,
            GLOBALBUFFEROUTPUT => \CLK_0_c_g\
        );

    \CLK_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2484\,
            DIN => \N__2483\,
            DOUT => \N__2482\,
            PACKAGEPIN => \CLK_wire\
        );

    \CLK_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__2484\,
            PADOUT => \N__2483\,
            PADIN => \N__2482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2473\,
            DIN => \N__2472\,
            DOUT => \N__2471\,
            PACKAGEPIN => \LED4_wire\
        );

    \LED4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2473\,
            PADOUT => \N__2472\,
            PADIN => \N__2471\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1212\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2464\,
            DIN => \N__2463\,
            DOUT => \N__2462\,
            PACKAGEPIN => \LED2_wire\
        );

    \LED2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2464\,
            PADOUT => \N__2463\,
            PADIN => \N__2462\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1284\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2455\,
            DIN => \N__2454\,
            DOUT => \N__2453\,
            PACKAGEPIN => \LED0_wire\
        );

    \LED0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2455\,
            PADOUT => \N__2454\,
            PADIN => \N__2453\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1326\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED6_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2446\,
            DIN => \N__2445\,
            DOUT => \N__2444\,
            PACKAGEPIN => \LED6_wire\
        );

    \LED6_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2446\,
            PADOUT => \N__2445\,
            PADIN => \N__2444\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1836\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2437\,
            DIN => \N__2436\,
            DOUT => \N__2435\,
            PACKAGEPIN => \LED3_wire\
        );

    \LED3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2437\,
            PADOUT => \N__2436\,
            PADIN => \N__2435\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1245\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED7_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2428\,
            DIN => \N__2427\,
            DOUT => \N__2426\,
            PACKAGEPIN => \LED7_wire\
        );

    \LED7_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2428\,
            PADOUT => \N__2427\,
            PADIN => \N__2426\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1740\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2419\,
            DIN => \N__2418\,
            DOUT => \N__2417\,
            PACKAGEPIN => \LED1_wire\
        );

    \LED1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2419\,
            PADOUT => \N__2418\,
            PADIN => \N__2417\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1977\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED5_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__2410\,
            DIN => \N__2409\,
            DOUT => \N__2408\,
            PACKAGEPIN => \LED5_wire\
        );

    \LED5_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__2410\,
            PADOUT => \N__2409\,
            PADIN => \N__2408\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__1176\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__2391\,
            I => \N__2387\
        );

    \I__522\ : InMux
    port map (
            O => \N__2390\,
            I => \N__2384\
        );

    \I__521\ : InMux
    port map (
            O => \N__2387\,
            I => \N__2381\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__2384\,
            I => \clk_divZ0Z_12\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__2381\,
            I => \clk_divZ0Z_12\
        );

    \I__518\ : InMux
    port map (
            O => \N__2376\,
            I => clk_div_1_cry_11
        );

    \I__517\ : CascadeMux
    port map (
            O => \N__2373\,
            I => \N__2369\
        );

    \I__516\ : InMux
    port map (
            O => \N__2372\,
            I => \N__2366\
        );

    \I__515\ : InMux
    port map (
            O => \N__2369\,
            I => \N__2363\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__2366\,
            I => \clk_divZ0Z_13\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__2363\,
            I => \clk_divZ0Z_13\
        );

    \I__512\ : InMux
    port map (
            O => \N__2358\,
            I => clk_div_1_cry_12
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__2355\,
            I => \N__2351\
        );

    \I__510\ : InMux
    port map (
            O => \N__2354\,
            I => \N__2348\
        );

    \I__509\ : InMux
    port map (
            O => \N__2351\,
            I => \N__2345\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__2348\,
            I => \clk_divZ0Z_14\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__2345\,
            I => \clk_divZ0Z_14\
        );

    \I__506\ : InMux
    port map (
            O => \N__2340\,
            I => clk_div_1_cry_13
        );

    \I__505\ : CascadeMux
    port map (
            O => \N__2337\,
            I => \N__2333\
        );

    \I__504\ : InMux
    port map (
            O => \N__2336\,
            I => \N__2330\
        );

    \I__503\ : InMux
    port map (
            O => \N__2333\,
            I => \N__2327\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__2330\,
            I => \clk_divZ0Z_15\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__2327\,
            I => \clk_divZ0Z_15\
        );

    \I__500\ : InMux
    port map (
            O => \N__2322\,
            I => clk_div_1_cry_14
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__2319\,
            I => \N__2315\
        );

    \I__498\ : InMux
    port map (
            O => \N__2318\,
            I => \N__2312\
        );

    \I__497\ : InMux
    port map (
            O => \N__2315\,
            I => \N__2309\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__2312\,
            I => \clk_divZ0Z_16\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__2309\,
            I => \clk_divZ0Z_16\
        );

    \I__494\ : InMux
    port map (
            O => \N__2304\,
            I => clk_div_1_cry_15
        );

    \I__493\ : CascadeMux
    port map (
            O => \N__2301\,
            I => \N__2297\
        );

    \I__492\ : InMux
    port map (
            O => \N__2300\,
            I => \N__2294\
        );

    \I__491\ : InMux
    port map (
            O => \N__2297\,
            I => \N__2291\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__2294\,
            I => \clk_divZ0Z_17\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__2291\,
            I => \clk_divZ0Z_17\
        );

    \I__488\ : InMux
    port map (
            O => \N__2286\,
            I => \bfn_2_11_0_\
        );

    \I__487\ : InMux
    port map (
            O => \N__2283\,
            I => clk_div_1_cry_17
        );

    \I__486\ : InMux
    port map (
            O => \N__2280\,
            I => \N__2276\
        );

    \I__485\ : InMux
    port map (
            O => \N__2279\,
            I => \N__2273\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__2276\,
            I => \clk_divZ0Z_18\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__2273\,
            I => \clk_divZ0Z_18\
        );

    \I__482\ : ClkMux
    port map (
            O => \N__2268\,
            I => \N__2244\
        );

    \I__481\ : ClkMux
    port map (
            O => \N__2267\,
            I => \N__2244\
        );

    \I__480\ : ClkMux
    port map (
            O => \N__2266\,
            I => \N__2244\
        );

    \I__479\ : ClkMux
    port map (
            O => \N__2265\,
            I => \N__2244\
        );

    \I__478\ : ClkMux
    port map (
            O => \N__2264\,
            I => \N__2244\
        );

    \I__477\ : ClkMux
    port map (
            O => \N__2263\,
            I => \N__2244\
        );

    \I__476\ : ClkMux
    port map (
            O => \N__2262\,
            I => \N__2244\
        );

    \I__475\ : ClkMux
    port map (
            O => \N__2261\,
            I => \N__2244\
        );

    \I__474\ : GlobalMux
    port map (
            O => \N__2244\,
            I => \N__2241\
        );

    \I__473\ : gio2CtrlBuf
    port map (
            O => \N__2241\,
            I => \CLK_0_c_g\
        );

    \I__472\ : InMux
    port map (
            O => \N__2238\,
            I => clk_div_1_cry_2
        );

    \I__471\ : CascadeMux
    port map (
            O => \N__2235\,
            I => \N__2231\
        );

    \I__470\ : InMux
    port map (
            O => \N__2234\,
            I => \N__2228\
        );

    \I__469\ : InMux
    port map (
            O => \N__2231\,
            I => \N__2225\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__2228\,
            I => \clk_divZ0Z_4\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__2225\,
            I => \clk_divZ0Z_4\
        );

    \I__466\ : InMux
    port map (
            O => \N__2220\,
            I => clk_div_1_cry_3
        );

    \I__465\ : CascadeMux
    port map (
            O => \N__2217\,
            I => \N__2213\
        );

    \I__464\ : InMux
    port map (
            O => \N__2216\,
            I => \N__2210\
        );

    \I__463\ : InMux
    port map (
            O => \N__2213\,
            I => \N__2207\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__2210\,
            I => \clk_divZ0Z_5\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__2207\,
            I => \clk_divZ0Z_5\
        );

    \I__460\ : InMux
    port map (
            O => \N__2202\,
            I => clk_div_1_cry_4
        );

    \I__459\ : CascadeMux
    port map (
            O => \N__2199\,
            I => \N__2195\
        );

    \I__458\ : InMux
    port map (
            O => \N__2198\,
            I => \N__2192\
        );

    \I__457\ : InMux
    port map (
            O => \N__2195\,
            I => \N__2189\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__2192\,
            I => \clk_divZ0Z_6\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__2189\,
            I => \clk_divZ0Z_6\
        );

    \I__454\ : InMux
    port map (
            O => \N__2184\,
            I => clk_div_1_cry_5
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__2181\,
            I => \N__2177\
        );

    \I__452\ : InMux
    port map (
            O => \N__2180\,
            I => \N__2174\
        );

    \I__451\ : InMux
    port map (
            O => \N__2177\,
            I => \N__2171\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__2174\,
            I => \clk_divZ0Z_7\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2171\,
            I => \clk_divZ0Z_7\
        );

    \I__448\ : InMux
    port map (
            O => \N__2166\,
            I => clk_div_1_cry_6
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__2163\,
            I => \N__2159\
        );

    \I__446\ : InMux
    port map (
            O => \N__2162\,
            I => \N__2156\
        );

    \I__445\ : InMux
    port map (
            O => \N__2159\,
            I => \N__2153\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2156\,
            I => \clk_divZ0Z_8\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__2153\,
            I => \clk_divZ0Z_8\
        );

    \I__442\ : InMux
    port map (
            O => \N__2148\,
            I => clk_div_1_cry_7
        );

    \I__441\ : CascadeMux
    port map (
            O => \N__2145\,
            I => \N__2141\
        );

    \I__440\ : InMux
    port map (
            O => \N__2144\,
            I => \N__2138\
        );

    \I__439\ : InMux
    port map (
            O => \N__2141\,
            I => \N__2135\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__2138\,
            I => \clk_divZ0Z_9\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__2135\,
            I => \clk_divZ0Z_9\
        );

    \I__436\ : InMux
    port map (
            O => \N__2130\,
            I => \bfn_2_10_0_\
        );

    \I__435\ : CascadeMux
    port map (
            O => \N__2127\,
            I => \N__2123\
        );

    \I__434\ : InMux
    port map (
            O => \N__2126\,
            I => \N__2120\
        );

    \I__433\ : InMux
    port map (
            O => \N__2123\,
            I => \N__2117\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__2120\,
            I => \clk_divZ0Z_10\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2117\,
            I => \clk_divZ0Z_10\
        );

    \I__430\ : InMux
    port map (
            O => \N__2112\,
            I => clk_div_1_cry_9
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__2109\,
            I => \N__2105\
        );

    \I__428\ : InMux
    port map (
            O => \N__2108\,
            I => \N__2102\
        );

    \I__427\ : InMux
    port map (
            O => \N__2105\,
            I => \N__2099\
        );

    \I__426\ : LocalMux
    port map (
            O => \N__2102\,
            I => \clk_divZ0Z_11\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2099\,
            I => \clk_divZ0Z_11\
        );

    \I__424\ : InMux
    port map (
            O => \N__2094\,
            I => clk_div_1_cry_10
        );

    \I__423\ : InMux
    port map (
            O => \N__2091\,
            I => \N__2086\
        );

    \I__422\ : InMux
    port map (
            O => \N__2090\,
            I => \N__2081\
        );

    \I__421\ : InMux
    port map (
            O => \N__2089\,
            I => \N__2081\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__2086\,
            I => \N__2076\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__2081\,
            I => \N__2076\
        );

    \I__418\ : Span4Mux_h
    port map (
            O => \N__2076\,
            I => \N__2072\
        );

    \I__417\ : InMux
    port map (
            O => \N__2075\,
            I => \N__2069\
        );

    \I__416\ : Odrv4
    port map (
            O => \N__2072\,
            I => clk_div_i_19
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2069\,
            I => clk_div_i_19
        );

    \I__414\ : InMux
    port map (
            O => \N__2064\,
            I => \N__2054\
        );

    \I__413\ : InMux
    port map (
            O => \N__2063\,
            I => \N__2047\
        );

    \I__412\ : InMux
    port map (
            O => \N__2062\,
            I => \N__2047\
        );

    \I__411\ : InMux
    port map (
            O => \N__2061\,
            I => \N__2047\
        );

    \I__410\ : InMux
    port map (
            O => \N__2060\,
            I => \N__2042\
        );

    \I__409\ : InMux
    port map (
            O => \N__2059\,
            I => \N__2042\
        );

    \I__408\ : InMux
    port map (
            O => \N__2058\,
            I => \N__2037\
        );

    \I__407\ : InMux
    port map (
            O => \N__2057\,
            I => \N__2037\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2054\,
            I => \cntrZ0Z_3\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2047\,
            I => \cntrZ0Z_3\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__2042\,
            I => \cntrZ0Z_3\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__2037\,
            I => \cntrZ0Z_3\
        );

    \I__402\ : CascadeMux
    port map (
            O => \N__2028\,
            I => \N__2024\
        );

    \I__401\ : InMux
    port map (
            O => \N__2027\,
            I => \N__2019\
        );

    \I__400\ : InMux
    port map (
            O => \N__2024\,
            I => \N__2016\
        );

    \I__399\ : InMux
    port map (
            O => \N__2023\,
            I => \N__2011\
        );

    \I__398\ : InMux
    port map (
            O => \N__2022\,
            I => \N__2011\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__2019\,
            I => \N_22\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__2016\,
            I => \N_22\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2011\,
            I => \N_22\
        );

    \I__394\ : InMux
    port map (
            O => \N__2004\,
            I => \N__2001\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__2001\,
            I => \N_21\
        );

    \I__392\ : InMux
    port map (
            O => \N__1998\,
            I => \N__1989\
        );

    \I__391\ : InMux
    port map (
            O => \N__1997\,
            I => \N__1989\
        );

    \I__390\ : InMux
    port map (
            O => \N__1996\,
            I => \N__1989\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__1989\,
            I => \N__1985\
        );

    \I__388\ : InMux
    port map (
            O => \N__1988\,
            I => \N__1982\
        );

    \I__387\ : Odrv4
    port map (
            O => \N__1985\,
            I => \N_19\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__1982\,
            I => \N_19\
        );

    \I__385\ : IoInMux
    port map (
            O => \N__1977\,
            I => \N__1973\
        );

    \I__384\ : CascadeMux
    port map (
            O => \N__1976\,
            I => \N__1970\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__1973\,
            I => \N__1967\
        );

    \I__382\ : InMux
    port map (
            O => \N__1970\,
            I => \N__1963\
        );

    \I__381\ : Span4Mux_s0_h
    port map (
            O => \N__1967\,
            I => \N__1960\
        );

    \I__380\ : InMux
    port map (
            O => \N__1966\,
            I => \N__1957\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__1963\,
            I => \N__1954\
        );

    \I__378\ : Odrv4
    port map (
            O => \N__1960\,
            I => \LED1_c\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__1957\,
            I => \LED1_c\
        );

    \I__376\ : Odrv4
    port map (
            O => \N__1954\,
            I => \LED1_c\
        );

    \I__375\ : InMux
    port map (
            O => \N__1947\,
            I => \N__1941\
        );

    \I__374\ : InMux
    port map (
            O => \N__1946\,
            I => \N__1941\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__1941\,
            I => \N_38\
        );

    \I__372\ : InMux
    port map (
            O => \N__1938\,
            I => \N__1935\
        );

    \I__371\ : LocalMux
    port map (
            O => \N__1935\,
            I => \BIT_47_1\
        );

    \I__370\ : InMux
    port map (
            O => \N__1932\,
            I => \N__1927\
        );

    \I__369\ : CascadeMux
    port map (
            O => \N__1931\,
            I => \N__1923\
        );

    \I__368\ : InMux
    port map (
            O => \N__1930\,
            I => \N__1919\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__1927\,
            I => \N__1916\
        );

    \I__366\ : InMux
    port map (
            O => \N__1926\,
            I => \N__1913\
        );

    \I__365\ : InMux
    port map (
            O => \N__1923\,
            I => \N__1908\
        );

    \I__364\ : InMux
    port map (
            O => \N__1922\,
            I => \N__1908\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__1919\,
            I => \cntrZ0Z_4\
        );

    \I__362\ : Odrv4
    port map (
            O => \N__1916\,
            I => \cntrZ0Z_4\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__1913\,
            I => \cntrZ0Z_4\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__1908\,
            I => \cntrZ0Z_4\
        );

    \I__359\ : InMux
    port map (
            O => \N__1899\,
            I => \N__1896\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__1896\,
            I => \N__1893\
        );

    \I__357\ : Odrv4
    port map (
            O => \N__1893\,
            I => g0_0
        );

    \I__356\ : CascadeMux
    port map (
            O => \N__1890\,
            I => \N__1887\
        );

    \I__355\ : InMux
    port map (
            O => \N__1887\,
            I => \N__1884\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__1884\,
            I => g0_4
        );

    \I__353\ : CascadeMux
    port map (
            O => \N__1881\,
            I => \N__1876\
        );

    \I__352\ : InMux
    port map (
            O => \N__1880\,
            I => \N__1872\
        );

    \I__351\ : InMux
    port map (
            O => \N__1879\,
            I => \N__1869\
        );

    \I__350\ : InMux
    port map (
            O => \N__1876\,
            I => \N__1866\
        );

    \I__349\ : InMux
    port map (
            O => \N__1875\,
            I => \N__1863\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__1872\,
            I => \N__1860\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__1869\,
            I => \N__1857\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__1866\,
            I => \N__1854\
        );

    \I__345\ : LocalMux
    port map (
            O => \N__1863\,
            I => \clk_div_RNIK8D95Z0Z_19\
        );

    \I__344\ : Odrv4
    port map (
            O => \N__1860\,
            I => \clk_div_RNIK8D95Z0Z_19\
        );

    \I__343\ : Odrv4
    port map (
            O => \N__1857\,
            I => \clk_div_RNIK8D95Z0Z_19\
        );

    \I__342\ : Odrv4
    port map (
            O => \N__1854\,
            I => \clk_div_RNIK8D95Z0Z_19\
        );

    \I__341\ : CascadeMux
    port map (
            O => \N__1845\,
            I => \cntr_RNIVLLQ5Z0Z_4_cascade_\
        );

    \I__340\ : InMux
    port map (
            O => \N__1842\,
            I => \N__1839\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__1839\,
            I => \BIT_47_6\
        );

    \I__338\ : IoInMux
    port map (
            O => \N__1836\,
            I => \N__1833\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__1833\,
            I => \N__1829\
        );

    \I__336\ : InMux
    port map (
            O => \N__1832\,
            I => \N__1825\
        );

    \I__335\ : Span4Mux_s3_v
    port map (
            O => \N__1829\,
            I => \N__1822\
        );

    \I__334\ : InMux
    port map (
            O => \N__1828\,
            I => \N__1819\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__1825\,
            I => \N__1816\
        );

    \I__332\ : Odrv4
    port map (
            O => \N__1822\,
            I => \LED6_c\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__1819\,
            I => \LED6_c\
        );

    \I__330\ : Odrv4
    port map (
            O => \N__1816\,
            I => \LED6_c\
        );

    \I__329\ : InMux
    port map (
            O => \N__1809\,
            I => \N__1797\
        );

    \I__328\ : InMux
    port map (
            O => \N__1808\,
            I => \N__1797\
        );

    \I__327\ : CEMux
    port map (
            O => \N__1807\,
            I => \N__1794\
        );

    \I__326\ : InMux
    port map (
            O => \N__1806\,
            I => \N__1783\
        );

    \I__325\ : InMux
    port map (
            O => \N__1805\,
            I => \N__1783\
        );

    \I__324\ : InMux
    port map (
            O => \N__1804\,
            I => \N__1783\
        );

    \I__323\ : InMux
    port map (
            O => \N__1803\,
            I => \N__1783\
        );

    \I__322\ : InMux
    port map (
            O => \N__1802\,
            I => \N__1783\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__1797\,
            I => \clk_div_RNIICCP5Z0Z_19\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__1794\,
            I => \clk_div_RNIICCP5Z0Z_19\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__1783\,
            I => \clk_div_RNIICCP5Z0Z_19\
        );

    \I__318\ : CascadeMux
    port map (
            O => \N__1776\,
            I => \N__1773\
        );

    \I__317\ : InMux
    port map (
            O => \N__1773\,
            I => \N__1770\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__1770\,
            I => \BIT_47_7\
        );

    \I__315\ : InMux
    port map (
            O => \N__1767\,
            I => \N__1758\
        );

    \I__314\ : InMux
    port map (
            O => \N__1766\,
            I => \N__1745\
        );

    \I__313\ : InMux
    port map (
            O => \N__1765\,
            I => \N__1745\
        );

    \I__312\ : InMux
    port map (
            O => \N__1764\,
            I => \N__1745\
        );

    \I__311\ : InMux
    port map (
            O => \N__1763\,
            I => \N__1745\
        );

    \I__310\ : InMux
    port map (
            O => \N__1762\,
            I => \N__1745\
        );

    \I__309\ : InMux
    port map (
            O => \N__1761\,
            I => \N__1745\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__1758\,
            I => \cntr_RNIVLLQ5Z0Z_4\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__1745\,
            I => \cntr_RNIVLLQ5Z0Z_4\
        );

    \I__306\ : IoInMux
    port map (
            O => \N__1740\,
            I => \N__1737\
        );

    \I__305\ : LocalMux
    port map (
            O => \N__1737\,
            I => \N__1733\
        );

    \I__304\ : CascadeMux
    port map (
            O => \N__1736\,
            I => \N__1730\
        );

    \I__303\ : IoSpan4Mux
    port map (
            O => \N__1733\,
            I => \N__1726\
        );

    \I__302\ : InMux
    port map (
            O => \N__1730\,
            I => \N__1723\
        );

    \I__301\ : InMux
    port map (
            O => \N__1729\,
            I => \N__1720\
        );

    \I__300\ : Span4Mux_s1_h
    port map (
            O => \N__1726\,
            I => \N__1715\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__1723\,
            I => \N__1715\
        );

    \I__298\ : LocalMux
    port map (
            O => \N__1720\,
            I => \LED7_c\
        );

    \I__297\ : Odrv4
    port map (
            O => \N__1715\,
            I => \LED7_c\
        );

    \I__296\ : SRMux
    port map (
            O => \N__1710\,
            I => \N__1706\
        );

    \I__295\ : SRMux
    port map (
            O => \N__1709\,
            I => \N__1703\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__1706\,
            I => \N__1700\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__1703\,
            I => \N__1697\
        );

    \I__292\ : Span4Mux_s2_h
    port map (
            O => \N__1700\,
            I => \N__1694\
        );

    \I__291\ : Odrv4
    port map (
            O => \N__1697\,
            I => \clk_div_RNI0HSQ5Z0Z_19\
        );

    \I__290\ : Odrv4
    port map (
            O => \N__1694\,
            I => \clk_div_RNI0HSQ5Z0Z_19\
        );

    \I__289\ : InMux
    port map (
            O => \N__1689\,
            I => \N__1685\
        );

    \I__288\ : InMux
    port map (
            O => \N__1688\,
            I => \N__1681\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__1685\,
            I => \N__1678\
        );

    \I__286\ : InMux
    port map (
            O => \N__1684\,
            I => \N__1675\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__1681\,
            I => \clk_divZ0Z_1\
        );

    \I__284\ : Odrv4
    port map (
            O => \N__1678\,
            I => \clk_divZ0Z_1\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__1675\,
            I => \clk_divZ0Z_1\
        );

    \I__282\ : CascadeMux
    port map (
            O => \N__1668\,
            I => \N__1665\
        );

    \I__281\ : InMux
    port map (
            O => \N__1665\,
            I => \N__1659\
        );

    \I__280\ : CascadeMux
    port map (
            O => \N__1664\,
            I => \N__1656\
        );

    \I__279\ : InMux
    port map (
            O => \N__1663\,
            I => \N__1651\
        );

    \I__278\ : InMux
    port map (
            O => \N__1662\,
            I => \N__1651\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__1659\,
            I => \N__1648\
        );

    \I__276\ : InMux
    port map (
            O => \N__1656\,
            I => \N__1645\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__1651\,
            I => \clk_divZ0Z_0\
        );

    \I__274\ : Odrv4
    port map (
            O => \N__1648\,
            I => \clk_divZ0Z_0\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__1645\,
            I => \clk_divZ0Z_0\
        );

    \I__272\ : CascadeMux
    port map (
            O => \N__1638\,
            I => \N__1634\
        );

    \I__271\ : InMux
    port map (
            O => \N__1637\,
            I => \N__1631\
        );

    \I__270\ : InMux
    port map (
            O => \N__1634\,
            I => \N__1628\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__1631\,
            I => \clk_divZ0Z_2\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__1628\,
            I => \clk_divZ0Z_2\
        );

    \I__267\ : InMux
    port map (
            O => \N__1623\,
            I => clk_div_1_cry_1
        );

    \I__266\ : CascadeMux
    port map (
            O => \N__1620\,
            I => \N__1616\
        );

    \I__265\ : InMux
    port map (
            O => \N__1619\,
            I => \N__1613\
        );

    \I__264\ : InMux
    port map (
            O => \N__1616\,
            I => \N__1610\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__1613\,
            I => \clk_divZ0Z_3\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__1610\,
            I => \clk_divZ0Z_3\
        );

    \I__261\ : InMux
    port map (
            O => \N__1605\,
            I => cntr_cry_3
        );

    \I__260\ : InMux
    port map (
            O => \N__1602\,
            I => cntr_cry_4
        );

    \I__259\ : InMux
    port map (
            O => \N__1599\,
            I => cntr_cry_5
        );

    \I__258\ : CascadeMux
    port map (
            O => \N__1596\,
            I => \N__1589\
        );

    \I__257\ : InMux
    port map (
            O => \N__1595\,
            I => \N__1584\
        );

    \I__256\ : InMux
    port map (
            O => \N__1594\,
            I => \N__1579\
        );

    \I__255\ : InMux
    port map (
            O => \N__1593\,
            I => \N__1579\
        );

    \I__254\ : InMux
    port map (
            O => \N__1592\,
            I => \N__1574\
        );

    \I__253\ : InMux
    port map (
            O => \N__1589\,
            I => \N__1574\
        );

    \I__252\ : InMux
    port map (
            O => \N__1588\,
            I => \N__1569\
        );

    \I__251\ : InMux
    port map (
            O => \N__1587\,
            I => \N__1569\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__1584\,
            I => \cntrZ0Z_6\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__1579\,
            I => \cntrZ0Z_6\
        );

    \I__248\ : LocalMux
    port map (
            O => \N__1574\,
            I => \cntrZ0Z_6\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__1569\,
            I => \cntrZ0Z_6\
        );

    \I__246\ : InMux
    port map (
            O => \N__1560\,
            I => \N__1557\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__1557\,
            I => \N__1553\
        );

    \I__244\ : InMux
    port map (
            O => \N__1556\,
            I => \N__1550\
        );

    \I__243\ : Odrv4
    port map (
            O => \N__1553\,
            I => \N_23\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__1550\,
            I => \N_23\
        );

    \I__241\ : InMux
    port map (
            O => \N__1545\,
            I => \N__1538\
        );

    \I__240\ : InMux
    port map (
            O => \N__1544\,
            I => \N__1535\
        );

    \I__239\ : InMux
    port map (
            O => \N__1543\,
            I => \N__1532\
        );

    \I__238\ : InMux
    port map (
            O => \N__1542\,
            I => \N__1527\
        );

    \I__237\ : InMux
    port map (
            O => \N__1541\,
            I => \N__1527\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__1538\,
            I => \cntrZ0Z_2\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__1535\,
            I => \cntrZ0Z_2\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__1532\,
            I => \cntrZ0Z_2\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__1527\,
            I => \cntrZ0Z_2\
        );

    \I__232\ : CascadeMux
    port map (
            O => \N__1518\,
            I => \N_21_cascade_\
        );

    \I__231\ : CascadeMux
    port map (
            O => \N__1515\,
            I => \N__1511\
        );

    \I__230\ : InMux
    port map (
            O => \N__1514\,
            I => \N__1502\
        );

    \I__229\ : InMux
    port map (
            O => \N__1511\,
            I => \N__1499\
        );

    \I__228\ : InMux
    port map (
            O => \N__1510\,
            I => \N__1494\
        );

    \I__227\ : InMux
    port map (
            O => \N__1509\,
            I => \N__1494\
        );

    \I__226\ : InMux
    port map (
            O => \N__1508\,
            I => \N__1489\
        );

    \I__225\ : InMux
    port map (
            O => \N__1507\,
            I => \N__1489\
        );

    \I__224\ : InMux
    port map (
            O => \N__1506\,
            I => \N__1484\
        );

    \I__223\ : InMux
    port map (
            O => \N__1505\,
            I => \N__1484\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__1502\,
            I => \cntrZ0Z_5\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__1499\,
            I => \cntrZ0Z_5\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__1494\,
            I => \cntrZ0Z_5\
        );

    \I__219\ : LocalMux
    port map (
            O => \N__1489\,
            I => \cntrZ0Z_5\
        );

    \I__218\ : LocalMux
    port map (
            O => \N__1484\,
            I => \cntrZ0Z_5\
        );

    \I__217\ : InMux
    port map (
            O => \N__1473\,
            I => \N__1466\
        );

    \I__216\ : InMux
    port map (
            O => \N__1472\,
            I => \N__1463\
        );

    \I__215\ : InMux
    port map (
            O => \N__1471\,
            I => \N__1458\
        );

    \I__214\ : InMux
    port map (
            O => \N__1470\,
            I => \N__1458\
        );

    \I__213\ : InMux
    port map (
            O => \N__1469\,
            I => \N__1455\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__1466\,
            I => \cntrZ0Z_0\
        );

    \I__211\ : LocalMux
    port map (
            O => \N__1463\,
            I => \cntrZ0Z_0\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__1458\,
            I => \cntrZ0Z_0\
        );

    \I__209\ : LocalMux
    port map (
            O => \N__1455\,
            I => \cntrZ0Z_0\
        );

    \I__208\ : CascadeMux
    port map (
            O => \N__1446\,
            I => \BIT_47_i_o3_0_0_4_cascade_\
        );

    \I__207\ : CascadeMux
    port map (
            O => \N__1443\,
            I => \N__1437\
        );

    \I__206\ : InMux
    port map (
            O => \N__1442\,
            I => \N__1434\
        );

    \I__205\ : InMux
    port map (
            O => \N__1441\,
            I => \N__1427\
        );

    \I__204\ : InMux
    port map (
            O => \N__1440\,
            I => \N__1427\
        );

    \I__203\ : InMux
    port map (
            O => \N__1437\,
            I => \N__1427\
        );

    \I__202\ : LocalMux
    port map (
            O => \N__1434\,
            I => \N_27\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__1427\,
            I => \N_27\
        );

    \I__200\ : InMux
    port map (
            O => \N__1422\,
            I => \N__1410\
        );

    \I__199\ : InMux
    port map (
            O => \N__1421\,
            I => \N__1410\
        );

    \I__198\ : InMux
    port map (
            O => \N__1420\,
            I => \N__1410\
        );

    \I__197\ : InMux
    port map (
            O => \N__1419\,
            I => \N__1410\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__1410\,
            I => \N_45\
        );

    \I__195\ : InMux
    port map (
            O => \N__1407\,
            I => \N__1402\
        );

    \I__194\ : InMux
    port map (
            O => \N__1406\,
            I => \N__1399\
        );

    \I__193\ : InMux
    port map (
            O => \N__1405\,
            I => \N__1396\
        );

    \I__192\ : LocalMux
    port map (
            O => \N__1402\,
            I => \N_17\
        );

    \I__191\ : LocalMux
    port map (
            O => \N__1399\,
            I => \N_17\
        );

    \I__190\ : LocalMux
    port map (
            O => \N__1396\,
            I => \N_17\
        );

    \I__189\ : CascadeMux
    port map (
            O => \N__1389\,
            I => \N_45_cascade_\
        );

    \I__188\ : CascadeMux
    port map (
            O => \N__1386\,
            I => \N__1383\
        );

    \I__187\ : InMux
    port map (
            O => \N__1383\,
            I => \N__1377\
        );

    \I__186\ : InMux
    port map (
            O => \N__1382\,
            I => \N__1377\
        );

    \I__185\ : LocalMux
    port map (
            O => \N__1377\,
            I => \N_30\
        );

    \I__184\ : InMux
    port map (
            O => \N__1374\,
            I => \bfn_2_6_0_\
        );

    \I__183\ : InMux
    port map (
            O => \N__1371\,
            I => \N__1364\
        );

    \I__182\ : InMux
    port map (
            O => \N__1370\,
            I => \N__1361\
        );

    \I__181\ : InMux
    port map (
            O => \N__1369\,
            I => \N__1356\
        );

    \I__180\ : InMux
    port map (
            O => \N__1368\,
            I => \N__1356\
        );

    \I__179\ : InMux
    port map (
            O => \N__1367\,
            I => \N__1353\
        );

    \I__178\ : LocalMux
    port map (
            O => \N__1364\,
            I => \cntrZ0Z_1\
        );

    \I__177\ : LocalMux
    port map (
            O => \N__1361\,
            I => \cntrZ0Z_1\
        );

    \I__176\ : LocalMux
    port map (
            O => \N__1356\,
            I => \cntrZ0Z_1\
        );

    \I__175\ : LocalMux
    port map (
            O => \N__1353\,
            I => \cntrZ0Z_1\
        );

    \I__174\ : InMux
    port map (
            O => \N__1344\,
            I => cntr_cry_0
        );

    \I__173\ : InMux
    port map (
            O => \N__1341\,
            I => cntr_cry_1
        );

    \I__172\ : InMux
    port map (
            O => \N__1338\,
            I => cntr_cry_2
        );

    \I__171\ : InMux
    port map (
            O => \N__1335\,
            I => clk_div_2_cry_18
        );

    \I__170\ : InMux
    port map (
            O => \N__1332\,
            I => \N__1329\
        );

    \I__169\ : LocalMux
    port map (
            O => \N__1329\,
            I => \BIT_47_0\
        );

    \I__168\ : IoInMux
    port map (
            O => \N__1326\,
            I => \N__1323\
        );

    \I__167\ : LocalMux
    port map (
            O => \N__1323\,
            I => \N__1320\
        );

    \I__166\ : Span4Mux_s2_v
    port map (
            O => \N__1320\,
            I => \N__1317\
        );

    \I__165\ : Span4Mux_v
    port map (
            O => \N__1317\,
            I => \N__1313\
        );

    \I__164\ : CascadeMux
    port map (
            O => \N__1316\,
            I => \N__1310\
        );

    \I__163\ : Span4Mux_h
    port map (
            O => \N__1313\,
            I => \N__1306\
        );

    \I__162\ : InMux
    port map (
            O => \N__1310\,
            I => \N__1303\
        );

    \I__161\ : InMux
    port map (
            O => \N__1309\,
            I => \N__1300\
        );

    \I__160\ : Odrv4
    port map (
            O => \N__1306\,
            I => \LED0_c\
        );

    \I__159\ : LocalMux
    port map (
            O => \N__1303\,
            I => \LED0_c\
        );

    \I__158\ : LocalMux
    port map (
            O => \N__1300\,
            I => \LED0_c\
        );

    \I__157\ : CascadeMux
    port map (
            O => \N__1293\,
            I => \clk_div_RNIICCP5Z0Z_19_cascade_\
        );

    \I__156\ : InMux
    port map (
            O => \N__1290\,
            I => \N__1287\
        );

    \I__155\ : LocalMux
    port map (
            O => \N__1287\,
            I => \N_12_i\
        );

    \I__154\ : IoInMux
    port map (
            O => \N__1284\,
            I => \N__1281\
        );

    \I__153\ : LocalMux
    port map (
            O => \N__1281\,
            I => \N__1277\
        );

    \I__152\ : CascadeMux
    port map (
            O => \N__1280\,
            I => \N__1274\
        );

    \I__151\ : Span4Mux_s2_v
    port map (
            O => \N__1277\,
            I => \N__1270\
        );

    \I__150\ : InMux
    port map (
            O => \N__1274\,
            I => \N__1267\
        );

    \I__149\ : InMux
    port map (
            O => \N__1273\,
            I => \N__1264\
        );

    \I__148\ : Span4Mux_h
    port map (
            O => \N__1270\,
            I => \N__1261\
        );

    \I__147\ : LocalMux
    port map (
            O => \N__1267\,
            I => \N__1256\
        );

    \I__146\ : LocalMux
    port map (
            O => \N__1264\,
            I => \N__1256\
        );

    \I__145\ : Odrv4
    port map (
            O => \N__1261\,
            I => \LED2_c\
        );

    \I__144\ : Odrv4
    port map (
            O => \N__1256\,
            I => \LED2_c\
        );

    \I__143\ : InMux
    port map (
            O => \N__1251\,
            I => \N__1248\
        );

    \I__142\ : LocalMux
    port map (
            O => \N__1248\,
            I => \N_14_i\
        );

    \I__141\ : IoInMux
    port map (
            O => \N__1245\,
            I => \N__1242\
        );

    \I__140\ : LocalMux
    port map (
            O => \N__1242\,
            I => \N__1238\
        );

    \I__139\ : CascadeMux
    port map (
            O => \N__1241\,
            I => \N__1235\
        );

    \I__138\ : IoSpan4Mux
    port map (
            O => \N__1238\,
            I => \N__1231\
        );

    \I__137\ : InMux
    port map (
            O => \N__1235\,
            I => \N__1228\
        );

    \I__136\ : InMux
    port map (
            O => \N__1234\,
            I => \N__1225\
        );

    \I__135\ : Odrv4
    port map (
            O => \N__1231\,
            I => \LED3_c\
        );

    \I__134\ : LocalMux
    port map (
            O => \N__1228\,
            I => \LED3_c\
        );

    \I__133\ : LocalMux
    port map (
            O => \N__1225\,
            I => \LED3_c\
        );

    \I__132\ : InMux
    port map (
            O => \N__1218\,
            I => \N__1215\
        );

    \I__131\ : LocalMux
    port map (
            O => \N__1215\,
            I => \N_6_i\
        );

    \I__130\ : IoInMux
    port map (
            O => \N__1212\,
            I => \N__1209\
        );

    \I__129\ : LocalMux
    port map (
            O => \N__1209\,
            I => \N__1206\
        );

    \I__128\ : Span4Mux_s2_v
    port map (
            O => \N__1206\,
            I => \N__1202\
        );

    \I__127\ : CascadeMux
    port map (
            O => \N__1205\,
            I => \N__1199\
        );

    \I__126\ : Span4Mux_v
    port map (
            O => \N__1202\,
            I => \N__1195\
        );

    \I__125\ : InMux
    port map (
            O => \N__1199\,
            I => \N__1192\
        );

    \I__124\ : InMux
    port map (
            O => \N__1198\,
            I => \N__1189\
        );

    \I__123\ : Odrv4
    port map (
            O => \N__1195\,
            I => \LED4_c\
        );

    \I__122\ : LocalMux
    port map (
            O => \N__1192\,
            I => \LED4_c\
        );

    \I__121\ : LocalMux
    port map (
            O => \N__1189\,
            I => \LED4_c\
        );

    \I__120\ : InMux
    port map (
            O => \N__1182\,
            I => \N__1179\
        );

    \I__119\ : LocalMux
    port map (
            O => \N__1179\,
            I => \N_8_i\
        );

    \I__118\ : IoInMux
    port map (
            O => \N__1176\,
            I => \N__1172\
        );

    \I__117\ : CascadeMux
    port map (
            O => \N__1175\,
            I => \N__1169\
        );

    \I__116\ : LocalMux
    port map (
            O => \N__1172\,
            I => \N__1165\
        );

    \I__115\ : InMux
    port map (
            O => \N__1169\,
            I => \N__1162\
        );

    \I__114\ : InMux
    port map (
            O => \N__1168\,
            I => \N__1159\
        );

    \I__113\ : Span4Mux_s0_h
    port map (
            O => \N__1165\,
            I => \N__1152\
        );

    \I__112\ : LocalMux
    port map (
            O => \N__1162\,
            I => \N__1152\
        );

    \I__111\ : LocalMux
    port map (
            O => \N__1159\,
            I => \N__1152\
        );

    \I__110\ : Odrv4
    port map (
            O => \N__1152\,
            I => \LED5_c\
        );

    \I__109\ : CascadeMux
    port map (
            O => \N__1149\,
            I => \N_17_cascade_\
        );

    \I__108\ : CascadeMux
    port map (
            O => \N__1146\,
            I => \N_22_cascade_\
        );

    \I__107\ : CascadeMux
    port map (
            O => \N__1143\,
            I => \N__1140\
        );

    \I__106\ : InMux
    port map (
            O => \N__1140\,
            I => \N__1137\
        );

    \I__105\ : LocalMux
    port map (
            O => \N__1137\,
            I => \BIT_47_0_a3_0_1_6\
        );

    \I__104\ : CascadeMux
    port map (
            O => \N__1134\,
            I => \N__1131\
        );

    \I__103\ : InMux
    port map (
            O => \N__1131\,
            I => \N__1125\
        );

    \I__102\ : InMux
    port map (
            O => \N__1130\,
            I => \N__1125\
        );

    \I__101\ : LocalMux
    port map (
            O => \N__1125\,
            I => \N__1122\
        );

    \I__100\ : Odrv4
    port map (
            O => \N__1122\,
            I => \N_31\
        );

    \I__99\ : CascadeMux
    port map (
            O => \N__1119\,
            I => \BIT_47_0_a3_0_1_6_cascade_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_8_0_\
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => clk_div_2_cry_8,
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => clk_div_2_cry_16,
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => clk_div_1_cry_8,
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => clk_div_1_cry_16,
            carryinitout => \bfn_2_11_0_\
        );

    \IN_MUX_bfv_2_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_6_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \cntr_RNI1FK_0_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__1368\,
            in1 => \N__1470\,
            in2 => \_gnd_net_\,
            in3 => \N__2059\,
            lcout => \BIT_47_0_a3_0_1_6\,
            ltout => \BIT_47_0_a3_0_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_RNI9VF1_6_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000100010"
        )
    port map (
            in0 => \N__1592\,
            in1 => \N__1405\,
            in2 => \N__1119\,
            in3 => \N__1510\,
            lcout => \N_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_RNI3ND_2_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2060\,
            in2 => \_gnd_net_\,
            in3 => \N__1543\,
            lcout => \N_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_RNI8GR_0_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__1471\,
            in1 => \N__1509\,
            in2 => \N__1596\,
            in3 => \N__1369\,
            lcout => \N_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_RNIVID_0_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1469\,
            in2 => \_gnd_net_\,
            in3 => \N__1367\,
            lcout => \N_17\,
            ltout => \N_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_RNIC891_6_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__1587\,
            in1 => \N__1505\,
            in2 => \N__1149\,
            in3 => \N__1419\,
            lcout => \N_22\,
            ltout => \N_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \BIT_RNO_0_3_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011000000"
        )
    port map (
            in0 => \N__1234\,
            in1 => \N__1442\,
            in2 => \N__1146\,
            in3 => \N__1382\,
            lcout => \N_14_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_RNIE4G1_0_6_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__1588\,
            in1 => \N__1506\,
            in2 => \N__1143\,
            in3 => \N__1420\,
            lcout => \N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \BIT_RNO_0_0_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010110011"
        )
    port map (
            in0 => \N__1309\,
            in1 => \N__1556\,
            in2 => \N__2028\,
            in3 => \N__1988\,
            lcout => \BIT_47_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \BIT_RNO_0_2_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000111111"
        )
    port map (
            in0 => \N__1273\,
            in1 => \N__1421\,
            in2 => \N__1134\,
            in3 => \N__1440\,
            lcout => \N_12_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \BIT_RNO_0_5_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000111"
        )
    port map (
            in0 => \N__1422\,
            in1 => \N__1130\,
            in2 => \N__1443\,
            in3 => \N__1168\,
            lcout => \N_8_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \BIT_RNO_0_4_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000000"
        )
    port map (
            in0 => \N__2027\,
            in1 => \N__1198\,
            in2 => \N__1386\,
            in3 => \N__1441\,
            lcout => \N_6_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \BIT_0_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011011100"
        )
    port map (
            in0 => \N__1804\,
            in1 => \N__1763\,
            in2 => \N__1316\,
            in3 => \N__1332\,
            lcout => \LED0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2262\,
            ce => 'H',
            sr => \N__1709\
        );

    \clk_div_RNIICCP5_19_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2091\,
            in2 => \_gnd_net_\,
            in3 => \N__1879\,
            lcout => \clk_div_RNIICCP5Z0Z_19\,
            ltout => \clk_div_RNIICCP5Z0Z_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \BIT_1_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101100"
        )
    port map (
            in0 => \N__1938\,
            in1 => \N__1966\,
            in2 => \N__1293\,
            in3 => \N__1764\,
            lcout => \LED1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2262\,
            ce => 'H',
            sr => \N__1709\
        );

    \BIT_2_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111010111010"
        )
    port map (
            in0 => \N__1761\,
            in1 => \N__1802\,
            in2 => \N__1280\,
            in3 => \N__1290\,
            lcout => \LED2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2262\,
            ce => 'H',
            sr => \N__1709\
        );

    \BIT_3_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011011100"
        )
    port map (
            in0 => \N__1805\,
            in1 => \N__1765\,
            in2 => \N__1241\,
            in3 => \N__1251\,
            lcout => \LED3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2262\,
            ce => 'H',
            sr => \N__1709\
        );

    \BIT_4_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111010111010"
        )
    port map (
            in0 => \N__1762\,
            in1 => \N__1803\,
            in2 => \N__1205\,
            in3 => \N__1218\,
            lcout => \LED4_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2262\,
            ce => 'H',
            sr => \N__1709\
        );

    \BIT_5_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011011100"
        )
    port map (
            in0 => \N__1806\,
            in1 => \N__1766\,
            in2 => \N__1175\,
            in3 => \N__1182\,
            lcout => \LED5_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2262\,
            ce => 'H',
            sr => \N__1709\
        );

    \clk_div_RNI91U1_1_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1684\,
            in2 => \N__1664\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_8_0_\,
            carryout => clk_div_2_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIF3T2_2_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1638\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_1,
            carryout => clk_div_2_cry_2,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIM6S3_3_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__1620\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_2,
            carryout => clk_div_2_cry_3,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIUAR4_4_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2235\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_3,
            carryout => clk_div_2_cry_4,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNI7GQ5_5_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2217\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_4,
            carryout => clk_div_2_cry_5,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIHMP6_6_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2199\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_5,
            carryout => clk_div_2_cry_6,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNISTO7_7_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2181\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_6,
            carryout => clk_div_2_cry_7,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNI86O8_8_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2163\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_7,
            carryout => clk_div_2_cry_8,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNILFN9_9_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2145\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => clk_div_2_cry_9,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIAAMP_10_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2127\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_9,
            carryout => clk_div_2_cry_10,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNI06L91_11_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2109\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_10,
            carryout => clk_div_2_cry_11,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIN2KP1_12_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2391\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_11,
            carryout => clk_div_2_cry_12,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIF0J92_13_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2373\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_12,
            carryout => clk_div_2_cry_13,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNI8VHP2_14_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2355\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_13,
            carryout => clk_div_2_cry_14,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNI2VG93_15_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2337\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_14,
            carryout => clk_div_2_cry_15,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNITVFP3_16_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2319\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_15,
            carryout => clk_div_2_cry_16,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIP1F94_17_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2301\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => clk_div_2_cry_17,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIM4EP4_18_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2279\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => clk_div_2_cry_17,
            carryout => clk_div_2_cry_18,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNIK8D95_19_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2075\,
            in2 => \_gnd_net_\,
            in3 => \N__1335\,
            lcout => \clk_div_RNIK8D95Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_19_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1875\,
            lcout => clk_div_i_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2263\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_RNI6KK_2_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111111"
        )
    port map (
            in0 => \N__1542\,
            in1 => \_gnd_net_\,
            in2 => \N__1931\,
            in3 => \N__2057\,
            lcout => OPEN,
            ltout => \BIT_47_i_o3_0_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_RNIE4G1_6_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__1594\,
            in1 => \N__1507\,
            in2 => \N__1446\,
            in3 => \N__1407\,
            lcout => \N_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_RNI4OD_2_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1541\,
            in2 => \_gnd_net_\,
            in3 => \N__1922\,
            lcout => \N_45\,
            ltout => \N_45_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_RNI9591_3_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__1508\,
            in1 => \N__1406\,
            in2 => \N__1389\,
            in3 => \N__2058\,
            lcout => \N_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_RNI5PD_1_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1593\,
            in2 => \_gnd_net_\,
            in3 => \N__1370\,
            lcout => g0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_0_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1473\,
            in2 => \_gnd_net_\,
            in3 => \N__1374\,
            lcout => \cntrZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_2_6_0_\,
            carryout => cntr_cry_0,
            clk => \N__2267\,
            ce => \N__1807\,
            sr => \_gnd_net_\
        );

    \cntr_1_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1371\,
            in2 => \_gnd_net_\,
            in3 => \N__1344\,
            lcout => \cntrZ0Z_1\,
            ltout => OPEN,
            carryin => cntr_cry_0,
            carryout => cntr_cry_1,
            clk => \N__2267\,
            ce => \N__1807\,
            sr => \_gnd_net_\
        );

    \cntr_2_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1545\,
            in2 => \_gnd_net_\,
            in3 => \N__1341\,
            lcout => \cntrZ0Z_2\,
            ltout => OPEN,
            carryin => cntr_cry_1,
            carryout => cntr_cry_2,
            clk => \N__2267\,
            ce => \N__1807\,
            sr => \_gnd_net_\
        );

    \cntr_3_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2064\,
            in2 => \_gnd_net_\,
            in3 => \N__1338\,
            lcout => \cntrZ0Z_3\,
            ltout => OPEN,
            carryin => cntr_cry_2,
            carryout => cntr_cry_3,
            clk => \N__2267\,
            ce => \N__1807\,
            sr => \_gnd_net_\
        );

    \cntr_4_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1930\,
            in2 => \_gnd_net_\,
            in3 => \N__1605\,
            lcout => \cntrZ0Z_4\,
            ltout => OPEN,
            carryin => cntr_cry_3,
            carryout => cntr_cry_4,
            clk => \N__2267\,
            ce => \N__1807\,
            sr => \_gnd_net_\
        );

    \cntr_5_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1514\,
            in2 => \_gnd_net_\,
            in3 => \N__1602\,
            lcout => \cntrZ0Z_5\,
            ltout => OPEN,
            carryin => cntr_cry_4,
            carryout => cntr_cry_5,
            clk => \N__2267\,
            ce => \N__1807\,
            sr => \_gnd_net_\
        );

    \cntr_6_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1595\,
            in2 => \_gnd_net_\,
            in3 => \N__1599\,
            lcout => \cntrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2267\,
            ce => \N__1807\,
            sr => \_gnd_net_\
        );

    \BIT_RNO_0_7_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100010001"
        )
    port map (
            in0 => \N__1998\,
            in1 => \N__1560\,
            in2 => \N__1736\,
            in3 => \N__2023\,
            lcout => \BIT_47_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_1_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1662\,
            in2 => \_gnd_net_\,
            in3 => \N__1688\,
            lcout => \clk_divZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_RNI6KK_0_2_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__1926\,
            in1 => \N__2061\,
            in2 => \_gnd_net_\,
            in3 => \N__1544\,
            lcout => \N_21\,
            ltout => \N_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \BIT_RNO_0_6_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001010"
        )
    port map (
            in0 => \N__1832\,
            in1 => \N__1997\,
            in2 => \N__1518\,
            in3 => \N__1947\,
            lcout => \BIT_47_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNI3NJG_19_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__2089\,
            in1 => \N__2062\,
            in2 => \N__1515\,
            in3 => \N__1472\,
            lcout => g0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_0_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1663\,
            lcout => \clk_divZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2264\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_RNI0HSQ5_19_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__2090\,
            in1 => \N__2063\,
            in2 => \N__1881\,
            in3 => \N__2022\,
            lcout => \clk_div_RNI0HSQ5Z0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \BIT_RNO_0_1_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010000"
        )
    port map (
            in0 => \N__2004\,
            in1 => \N__1996\,
            in2 => \N__1976\,
            in3 => \N__1946\,
            lcout => \BIT_47_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cntr_RNIVLLQ5_4_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__1932\,
            in1 => \N__1899\,
            in2 => \N__1890\,
            in3 => \N__1880\,
            lcout => \cntr_RNIVLLQ5Z0Z_4\,
            ltout => \cntr_RNIVLLQ5Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \BIT_6_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011110100"
        )
    port map (
            in0 => \N__1808\,
            in1 => \N__1828\,
            in2 => \N__1845\,
            in3 => \N__1842\,
            lcout => \LED6_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2261\,
            ce => 'H',
            sr => \N__1710\
        );

    \BIT_7_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111100100"
        )
    port map (
            in0 => \N__1809\,
            in1 => \N__1729\,
            in2 => \N__1776\,
            in3 => \N__1767\,
            lcout => \LED7_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2261\,
            ce => 'H',
            sr => \N__1710\
        );

    \clk_div_1_cry_1_c_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1689\,
            in2 => \N__1668\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => clk_div_1_cry_1,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_2_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1637\,
            in2 => \_gnd_net_\,
            in3 => \N__1623\,
            lcout => \clk_divZ0Z_2\,
            ltout => OPEN,
            carryin => clk_div_1_cry_1,
            carryout => clk_div_1_cry_2,
            clk => \N__2265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_3_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1619\,
            in2 => \_gnd_net_\,
            in3 => \N__2238\,
            lcout => \clk_divZ0Z_3\,
            ltout => OPEN,
            carryin => clk_div_1_cry_2,
            carryout => clk_div_1_cry_3,
            clk => \N__2265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_4_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2234\,
            in2 => \_gnd_net_\,
            in3 => \N__2220\,
            lcout => \clk_divZ0Z_4\,
            ltout => OPEN,
            carryin => clk_div_1_cry_3,
            carryout => clk_div_1_cry_4,
            clk => \N__2265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_5_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2216\,
            in2 => \_gnd_net_\,
            in3 => \N__2202\,
            lcout => \clk_divZ0Z_5\,
            ltout => OPEN,
            carryin => clk_div_1_cry_4,
            carryout => clk_div_1_cry_5,
            clk => \N__2265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_6_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2198\,
            in2 => \_gnd_net_\,
            in3 => \N__2184\,
            lcout => \clk_divZ0Z_6\,
            ltout => OPEN,
            carryin => clk_div_1_cry_5,
            carryout => clk_div_1_cry_6,
            clk => \N__2265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_7_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2180\,
            in2 => \_gnd_net_\,
            in3 => \N__2166\,
            lcout => \clk_divZ0Z_7\,
            ltout => OPEN,
            carryin => clk_div_1_cry_6,
            carryout => clk_div_1_cry_7,
            clk => \N__2265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_8_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2162\,
            in2 => \_gnd_net_\,
            in3 => \N__2148\,
            lcout => \clk_divZ0Z_8\,
            ltout => OPEN,
            carryin => clk_div_1_cry_7,
            carryout => clk_div_1_cry_8,
            clk => \N__2265\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_9_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2144\,
            in2 => \_gnd_net_\,
            in3 => \N__2130\,
            lcout => \clk_divZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => clk_div_1_cry_9,
            clk => \N__2266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_10_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2126\,
            in2 => \_gnd_net_\,
            in3 => \N__2112\,
            lcout => \clk_divZ0Z_10\,
            ltout => OPEN,
            carryin => clk_div_1_cry_9,
            carryout => clk_div_1_cry_10,
            clk => \N__2266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_11_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2108\,
            in2 => \_gnd_net_\,
            in3 => \N__2094\,
            lcout => \clk_divZ0Z_11\,
            ltout => OPEN,
            carryin => clk_div_1_cry_10,
            carryout => clk_div_1_cry_11,
            clk => \N__2266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_12_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2390\,
            in2 => \_gnd_net_\,
            in3 => \N__2376\,
            lcout => \clk_divZ0Z_12\,
            ltout => OPEN,
            carryin => clk_div_1_cry_11,
            carryout => clk_div_1_cry_12,
            clk => \N__2266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_13_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2372\,
            in2 => \_gnd_net_\,
            in3 => \N__2358\,
            lcout => \clk_divZ0Z_13\,
            ltout => OPEN,
            carryin => clk_div_1_cry_12,
            carryout => clk_div_1_cry_13,
            clk => \N__2266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_14_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2354\,
            in2 => \_gnd_net_\,
            in3 => \N__2340\,
            lcout => \clk_divZ0Z_14\,
            ltout => OPEN,
            carryin => clk_div_1_cry_13,
            carryout => clk_div_1_cry_14,
            clk => \N__2266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_15_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2336\,
            in2 => \_gnd_net_\,
            in3 => \N__2322\,
            lcout => \clk_divZ0Z_15\,
            ltout => OPEN,
            carryin => clk_div_1_cry_14,
            carryout => clk_div_1_cry_15,
            clk => \N__2266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_16_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2318\,
            in2 => \_gnd_net_\,
            in3 => \N__2304\,
            lcout => \clk_divZ0Z_16\,
            ltout => OPEN,
            carryin => clk_div_1_cry_15,
            carryout => clk_div_1_cry_16,
            clk => \N__2266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_17_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2300\,
            in2 => \_gnd_net_\,
            in3 => \N__2286\,
            lcout => \clk_divZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_2_11_0_\,
            carryout => clk_div_1_cry_17,
            clk => \N__2268\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_div_18_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2280\,
            in2 => \_gnd_net_\,
            in3 => \N__2283\,
            lcout => \clk_divZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__2268\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
